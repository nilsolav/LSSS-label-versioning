netcdf mask {
	:date_created = "20200811T114628";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200811T114628";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 41;
			channels = 6;
			categories = 246;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  63.1, 14.0, 13.9, 61.2, 55.5, 60.3, 62.7, 64.2, 65.3, 64.1, 68.2, 32.7, 31.9, 65.3, 52.3, 53.9, 54.1, 62.8, 52.5, 52.9, 56.9, 54.7, 51.0, 55.3, 57.4, 49.6, 58.5, 55.5, 60.5, 68.6, 68.0, 60.4, 64.8, 61.4, 62.3, 11.2, 10.9,  9.8, 11.6, 61.2, 64.2;
			max_depth =  64.4, 26.9, 23.9, 65.0, 61.4, 62.3, 65.7, 65.8, 66.7, 65.8, 69.2, 35.8, 34.0, 72.3, 61.7, 66.7, 58.6, 68.4, 60.6, 54.0, 60.3, 57.8, 62.4, 64.7, 62.2, 57.2, 64.1, 61.8, 67.8, 69.7, 69.7, 63.1, 67.3, 63.9, 64.9, 31.3, 31.8, 31.9, 34.4, 63.2, 65.7;
			start_time = 128874388596773248, 128874400233209600, 128874400761334528, 128874398341334528, 128874401549303168, 128874402789303296, 128874402801334528, 128874395088804480, 128874391672867072, 128874392076773248, 128874393788804608, 128874397881334528, 128874395220835840, 128874406385240704, 128874408653209600, 128874409037272064, 128874409289303296, 128874409405240704, 128874409773209472, 128874409837272064, 128874410841334400, 128874410957271936, 128874412153209472, 128874412605240832, 128874414613209472, 128874415501334528, 128874416701334400, 128874417641334528, 128874420469303296, 128874416169303296, 128874421789303296, 128874428217271936, 128874422545240832, 128874427081334528, 128874430521334528, 128874425541334528, 128874425693209472, 128874430621334528, 128874432065240704, 128874423169303168, 128874423381334400;
			end_time = 128874388620835840, 128874400465240832, 128874401045240704, 128874398365240832, 128874401573209472, 128874402805240704, 128874402829303296, 128874395112866944, 128874391696773248, 128874392092867072, 128874393808804480, 128874397901334400, 128874395236773248, 128874406449303296, 128874408741334528, 128874409221334528, 128874409353209472, 128874409449303168, 128874409833209472, 128874409853209472, 128874410861334528, 128874410989303296, 128874412261334528, 128874412665240832, 128874414661334400, 128874415585240704, 128874416733209472, 128874417693209472, 128874420521334400, 128874416197272064, 128874421833209472, 128874428253209472, 128874422581334528, 128874427117272064, 128874430549303168, 128874425677271936, 128874426753209472, 128874430841334528, 128874432413209472, 128874423193209472, 128874423417271936;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21","Layer22","Layer23","Layer24","Layer25","Layer26","Layer27","Layer28","Layer29","Layer30","Layer31","Layer32","Layer33","Layer34","Layer35","Layer36","Layer37","Layer38","Layer39","Layer40","Layer41";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63;
			mask_times = {1.288743885967732e+17, 1.288743886008357e+17, 1.288743886048983e+17, 1.288743886088045e+17, 1.288743886128671e+17, 1.288743886167732e+17, 1.288743886208358e+17},
			             {1.288744002332096e+17, 1.288744002372719e+17, 1.288744002413345e+17, 1.288744002452407e+17, 1.288744002493032e+17, 1.288744002532095e+17, 1.288744002572719e+17, 1.288744002613345e+17, 1.288744002652407e+17, 1.288744002693033e+17, 1.288744002732095e+17, 1.288744002772719e+17, 1.288744002813345e+17, 1.288744002852407e+17, 1.288744002893032e+17, 1.288744002932095e+17, 1.288744002972719e+17, 1.288744003013345e+17, 1.288744003052407e+17, 1.288744003093033e+17, 1.288744003132095e+17, 1.288744003172721e+17, 1.288744003213345e+17, 1.288744003252407e+17, 1.288744003293033e+17, 1.288744003332095e+17, 1.288744003372719e+17, 1.288744003413345e+17, 1.288744003452407e+17, 1.288744003532095e+17, 1.288744003572721e+17, 1.288744003613345e+17, 1.288744003652407e+17, 1.288744003693033e+17, 1.288744003732095e+17, 1.288744003772721e+17, 1.288744003813345e+17, 1.288744003852407e+17, 1.288744003893033e+17, 1.288744003932095e+17, 1.288744003972721e+17, 1.288744004013344e+17, 1.288744004052408e+17, 1.288744004093033e+17, 1.288744004132095e+17, 1.288744004172721e+17, 1.288744004213344e+17, 1.288744004252407e+17, 1.288744004293032e+17, 1.288744004332095e+17, 1.288744004452408e+17, 1.288744004532096e+17, 1.288744004572719e+17, 1.288744004613344e+17, 1.288744004652408e+17},
			             {1.288744007613345e+17, 1.288744007652407e+17, 1.288744007693032e+17, 1.288744007732095e+17, 1.288744007772719e+17, 1.288744007813345e+17, 1.288744007852407e+17, 1.288744007893033e+17, 1.288744007932095e+17, 1.288744007972719e+17, 1.288744008013345e+17, 1.288744008052407e+17, 1.288744008093033e+17, 1.288744008132095e+17, 1.288744008172719e+17, 1.288744008213345e+17, 1.288744008252407e+17, 1.288744008293033e+17, 1.288744008332095e+17, 1.288744008372721e+17, 1.288744008413345e+17, 1.288744008452407e+17, 1.288744008493033e+17, 1.288744008532095e+17, 1.288744008572719e+17, 1.288744008613345e+17, 1.288744008652407e+17, 1.288744008693033e+17, 1.288744008732095e+17, 1.288744008772721e+17, 1.288744008813345e+17, 1.288744008852408e+17, 1.288744008893033e+17, 1.288744008932095e+17, 1.288744008972721e+17, 1.288744009013345e+17, 1.288744009052407e+17, 1.288744009093033e+17, 1.288744009132095e+17, 1.288744009172721e+17, 1.288744009213345e+17, 1.288744009252408e+17, 1.288744009293033e+17, 1.288744009332095e+17, 1.288744009372721e+17, 1.288744009413344e+17, 1.288744009452407e+17, 1.288744009493032e+17, 1.288744009532095e+17, 1.288744009572721e+17, 1.288744009613345e+17, 1.288744009652408e+17, 1.288744009693032e+17, 1.288744009732096e+17, 1.288744009772719e+17, 1.288744009813344e+17, 1.288744009852408e+17, 1.288744009893032e+17, 1.288744009932095e+17, 1.288744009972719e+17, 1.288744010013345e+17, 1.288744010052407e+17, 1.288744010093033e+17, 1.288744010132096e+17, 1.288744010172719e+17, 1.288744010213345e+17, 1.288744010252407e+17, 1.288744010293032e+17, 1.288744010332095e+17, 1.288744010372719e+17, 1.288744010413345e+17, 1.288744010452407e+17},
			             {1.288743983413345e+17, 1.288743983452407e+17, 1.288743983493033e+17, 1.288743983532095e+17, 1.288743983572721e+17, 1.288743983613344e+17, 1.288743983652408e+17},
			             {1.288744015493032e+17, 1.288744015532095e+17, 1.288744015572719e+17, 1.288744015613345e+17, 1.288744015652407e+17, 1.288744015693033e+17, 1.288744015732095e+17},
			             {1.288744027893033e+17, 1.288744027932096e+17, 1.288744027972719e+17, 1.288744028013345e+17, 1.288744028052407e+17},
			             {1.288744028013345e+17, 1.288744028052407e+17, 1.288744028093032e+17, 1.288744028132095e+17, 1.288744028172719e+17, 1.288744028213345e+17, 1.288744028252407e+17, 1.288744028293033e+17},
			             {1.288743950888045e+17, 1.288743950928669e+17, 1.288743950967732e+17, 1.288743951008357e+17, 1.288743951048983e+17, 1.288743951088045e+17, 1.288743951128669e+17},
			             {1.288743916728671e+17, 1.288743916767732e+17, 1.288743916808357e+17, 1.288743916848982e+17, 1.288743916888045e+17, 1.288743916928671e+17, 1.288743916967732e+17},
			             {1.288743920767732e+17, 1.288743920808357e+17, 1.288743920848983e+17, 1.288743920888045e+17, 1.288743920928671e+17},
			             {1.288743937888046e+17, 1.288743937928669e+17, 1.288743937967732e+17, 1.288743938008357e+17, 1.288743938048982e+17, 1.288743938088045e+17},
			             {1.288743978813345e+17, 1.288743978852408e+17, 1.288743978893032e+17, 1.288743978932095e+17, 1.288743978972721e+17, 1.288743979013344e+17},
			             {1.288743952208358e+17, 1.288743952248983e+17, 1.288743952288045e+17, 1.288743952328671e+17, 1.288743952367732e+17},
			             {1.288744063852407e+17, 1.288744063893033e+17, 1.288744063932095e+17, 1.288744063972719e+17, 1.288744064013345e+17, 1.288744064052407e+17, 1.288744064093033e+17, 1.288744064132095e+17, 1.288744064172719e+17, 1.288744064213345e+17, 1.288744064252407e+17, 1.288744064293033e+17, 1.288744064332095e+17, 1.288744064372721e+17, 1.288744064413345e+17, 1.288744064452407e+17, 1.288744064493033e+17},
			             {1.288744086532096e+17, 1.288744086572719e+17, 1.288744086613345e+17, 1.288744086652407e+17, 1.288744086693032e+17, 1.288744086732095e+17, 1.288744086772719e+17, 1.288744086813345e+17, 1.288744086852407e+17, 1.288744086893033e+17, 1.288744086932095e+17, 1.288744086972719e+17, 1.288744087013345e+17, 1.288744087052407e+17, 1.288744087093033e+17, 1.288744087132095e+17, 1.288744087172719e+17, 1.288744087213345e+17, 1.288744087252407e+17, 1.288744087293033e+17, 1.288744087332095e+17, 1.288744087372721e+17, 1.288744087413345e+17},
			             {1.288744090372721e+17, 1.288744090413345e+17, 1.288744090452408e+17, 1.288744090493033e+17, 1.288744090532095e+17, 1.288744090572721e+17, 1.288744090613344e+17, 1.288744090652407e+17, 1.288744090693033e+17, 1.288744090732095e+17, 1.288744090772721e+17, 1.288744090813345e+17, 1.288744090852408e+17, 1.288744090893032e+17, 1.288744090932095e+17, 1.288744090972721e+17, 1.288744091013344e+17, 1.288744091052408e+17, 1.288744091093032e+17, 1.288744091132095e+17, 1.288744091172719e+17, 1.288744091213345e+17, 1.288744091252408e+17, 1.288744091293032e+17, 1.288744091332096e+17, 1.288744091372719e+17, 1.288744091413345e+17, 1.288744091452407e+17, 1.288744091493032e+17, 1.288744091532095e+17, 1.288744091572719e+17, 1.288744091613345e+17, 1.288744091652407e+17, 1.288744091693033e+17, 1.288744091732095e+17, 1.288744091772719e+17, 1.288744091813345e+17, 1.288744091852407e+17, 1.288744091893032e+17, 1.288744091932095e+17, 1.288744091972719e+17, 1.288744092013345e+17, 1.288744092052407e+17, 1.288744092093033e+17, 1.288744092132095e+17, 1.288744092172721e+17, 1.288744092213345e+17},
			             {1.288744092893033e+17, 1.288744092932095e+17, 1.288744092972721e+17, 1.288744093013345e+17, 1.288744093052408e+17, 1.288744093093033e+17, 1.288744093132095e+17, 1.288744093172721e+17, 1.288744093213344e+17, 1.288744093252407e+17, 1.288744093293033e+17, 1.288744093332095e+17, 1.288744093372721e+17, 1.288744093413345e+17, 1.288744093452408e+17, 1.288744093493032e+17, 1.288744093532095e+17},
			             {1.288744094052407e+17, 1.288744094093032e+17, 1.288744094132095e+17, 1.288744094172719e+17, 1.288744094213345e+17, 1.288744094252407e+17, 1.288744094293033e+17, 1.288744094332095e+17, 1.288744094372719e+17, 1.288744094413345e+17, 1.288744094452407e+17, 1.288744094493032e+17},
			             {1.288744097732095e+17, 1.288744097772721e+17, 1.288744097813345e+17, 1.288744097852407e+17, 1.288744097893033e+17, 1.288744097932095e+17, 1.288744097972721e+17, 1.288744098013345e+17, 1.288744098052407e+17, 1.288744098093033e+17, 1.288744098132095e+17, 1.288744098172721e+17, 1.288744098213344e+17, 1.288744098252408e+17, 1.288744098293033e+17, 1.288744098332095e+17},
			             {1.288744098372721e+17, 1.288744098413344e+17, 1.288744098452407e+17, 1.288744098493032e+17, 1.288744098532095e+17},
			             {1.288744108413344e+17, 1.288744108452407e+17, 1.288744108493033e+17, 1.288744108532095e+17, 1.288744108572721e+17, 1.288744108613345e+17},
			             {1.288744109572719e+17, 1.288744109613345e+17, 1.288744109652407e+17, 1.288744109693032e+17, 1.288744109732095e+17, 1.288744109772719e+17, 1.288744109813345e+17, 1.288744109852407e+17, 1.288744109893033e+17},
			             {1.288744121532095e+17, 1.288744121572721e+17, 1.288744121613345e+17, 1.288744121652408e+17, 1.288744121693032e+17, 1.288744121732096e+17, 1.288744121772719e+17, 1.288744121813344e+17, 1.288744121852408e+17, 1.288744121893032e+17, 1.288744121932095e+17, 1.288744121972719e+17, 1.288744122013345e+17, 1.288744122052407e+17, 1.288744122093033e+17, 1.288744122132096e+17, 1.288744122172719e+17, 1.288744122213345e+17, 1.288744122252407e+17, 1.288744122293032e+17, 1.288744122332095e+17, 1.288744122372719e+17, 1.288744122413345e+17, 1.288744122452407e+17, 1.288744122493033e+17, 1.288744122532095e+17, 1.288744122572719e+17, 1.288744122613345e+17},
			             {1.288744126052408e+17, 1.288744126093033e+17, 1.288744126132095e+17, 1.288744126172721e+17, 1.288744126213344e+17, 1.288744126252407e+17, 1.288744126293033e+17, 1.288744126332095e+17, 1.288744126372721e+17, 1.288744126413345e+17, 1.288744126452408e+17, 1.288744126493032e+17, 1.288744126532095e+17, 1.288744126572721e+17, 1.288744126613344e+17, 1.288744126652408e+17},
			             {1.288744146132095e+17, 1.288744146172719e+17, 1.288744146213345e+17, 1.288744146252407e+17, 1.288744146293033e+17, 1.288744146332095e+17, 1.288744146372721e+17, 1.288744146413345e+17, 1.288744146452408e+17, 1.288744146493033e+17, 1.288744146532095e+17, 1.288744146572721e+17, 1.288744146613344e+17},
			             {1.288744155013345e+17, 1.288744155052408e+17, 1.288744155093032e+17, 1.288744155132096e+17, 1.288744155172719e+17, 1.288744155213345e+17, 1.288744155252407e+17, 1.288744155293032e+17, 1.288744155332095e+17, 1.288744155372719e+17, 1.288744155413345e+17, 1.288744155452407e+17, 1.288744155493033e+17, 1.288744155532095e+17, 1.288744155572719e+17, 1.288744155613345e+17, 1.288744155652407e+17, 1.288744155693032e+17, 1.288744155732095e+17, 1.288744155772719e+17, 1.288744155813345e+17, 1.288744155852407e+17},
			             {1.288744167013344e+17, 1.288744167052407e+17, 1.288744167093033e+17, 1.288744167132095e+17, 1.288744167172721e+17, 1.288744167213345e+17, 1.288744167252408e+17, 1.288744167293032e+17, 1.288744167332095e+17},
			             {1.288744176413345e+17, 1.288744176452407e+17, 1.288744176493033e+17, 1.288744176532095e+17, 1.288744176572719e+17, 1.288744176613345e+17, 1.288744176652407e+17, 1.288744176693033e+17, 1.288744176732095e+17, 1.288744176772721e+17, 1.288744176813345e+17, 1.288744176852407e+17, 1.288744176893033e+17, 1.288744176932095e+17},
			             {1.288744204693033e+17, 1.288744204732095e+17, 1.288744204772719e+17, 1.288744204813345e+17, 1.288744204852407e+17, 1.288744204893033e+17, 1.288744204932095e+17, 1.288744204972721e+17, 1.288744205013345e+17, 1.288744205052408e+17, 1.288744205093033e+17, 1.288744205132095e+17, 1.288744205172721e+17, 1.288744205213344e+17},
			             {1.288744161693033e+17, 1.288744161732095e+17, 1.288744161772721e+17, 1.288744161813345e+17, 1.288744161852407e+17, 1.288744161893033e+17, 1.288744161932095e+17, 1.288744161972721e+17},
			             {1.288744217893033e+17, 1.288744217932095e+17, 1.288744217972721e+17, 1.288744218013344e+17, 1.288744218052408e+17, 1.288744218093033e+17, 1.288744218132095e+17, 1.288744218172721e+17, 1.288744218213344e+17, 1.288744218252407e+17, 1.288744218293032e+17, 1.288744218332095e+17},
			             {1.288744282172719e+17, 1.288744282213345e+17, 1.288744282252408e+17, 1.288744282293032e+17, 1.288744282332096e+17, 1.288744282372719e+17, 1.288744282413345e+17, 1.288744282452407e+17, 1.288744282493032e+17, 1.288744282532095e+17},
			             {1.288744225452408e+17, 1.288744225493033e+17, 1.288744225532095e+17, 1.288744225572721e+17, 1.288744225613344e+17, 1.288744225652407e+17, 1.288744225693033e+17, 1.288744225732095e+17, 1.288744225772721e+17, 1.288744225813345e+17},
			             {1.288744270813345e+17, 1.288744270852407e+17, 1.288744270893033e+17, 1.288744270932095e+17, 1.288744270972721e+17, 1.288744271013345e+17, 1.288744271052407e+17, 1.288744271093033e+17, 1.288744271132095e+17, 1.288744271172721e+17},
			             {1.288744305213345e+17, 1.288744305252408e+17, 1.288744305293032e+17, 1.288744305332096e+17, 1.288744305372719e+17, 1.288744305413345e+17, 1.288744305452407e+17, 1.288744305493032e+17},
			             {1.288744255413345e+17, 1.288744255452407e+17, 1.288744255493033e+17, 1.288744255532095e+17, 1.288744255572719e+17, 1.288744255613345e+17, 1.288744255652407e+17, 1.288744255693033e+17, 1.288744255732095e+17, 1.288744255772721e+17, 1.288744255813345e+17, 1.288744255852407e+17, 1.288744255893033e+17, 1.288744255932095e+17, 1.288744255972721e+17, 1.288744256013345e+17, 1.288744256052407e+17, 1.288744256093033e+17, 1.288744256132095e+17, 1.288744256172721e+17, 1.288744256213344e+17, 1.288744256252408e+17, 1.288744256293033e+17, 1.288744256332095e+17, 1.288744256372721e+17, 1.288744256413344e+17, 1.288744256452407e+17, 1.288744256493032e+17, 1.288744256532095e+17, 1.288744256572721e+17, 1.288744256613345e+17, 1.288744256652408e+17, 1.288744256693032e+17, 1.288744256732096e+17, 1.288744256772719e+17},
			             {1.288744256932095e+17, 1.288744256972719e+17, 1.288744257013345e+17, 1.288744257052407e+17, 1.288744257093033e+17, 1.288744257132096e+17, 1.288744257172719e+17, 1.288744257213345e+17, 1.288744257252407e+17, 1.288744257293032e+17, 1.288744257332095e+17, 1.288744257372719e+17, 1.288744257413345e+17, 1.288744257452407e+17, 1.288744257493033e+17, 1.288744257532095e+17, 1.288744257572719e+17, 1.288744257613345e+17, 1.288744257652407e+17, 1.288744257693033e+17, 1.288744257732095e+17, 1.288744257772719e+17, 1.288744257813345e+17, 1.288744257852407e+17, 1.288744257893033e+17, 1.288744257932095e+17, 1.288744257972721e+17, 1.288744258013345e+17, 1.288744258052407e+17, 1.288744258093033e+17, 1.288744258132095e+17, 1.288744258172719e+17, 1.288744258213345e+17, 1.288744258252407e+17, 1.288744258293033e+17, 1.288744258332095e+17, 1.288744258372721e+17, 1.288744258413345e+17, 1.288744258452407e+17, 1.288744258493033e+17, 1.288744258532095e+17, 1.288744258572721e+17, 1.288744258613345e+17, 1.288744258652407e+17, 1.288744258693033e+17, 1.288744258732095e+17, 1.288744258772721e+17, 1.288744258813345e+17, 1.288744258852408e+17, 1.288744258893033e+17, 1.288744258932095e+17, 1.288744258972721e+17, 1.288744259013344e+17, 1.288744259052407e+17, 1.288744259093032e+17, 1.288744259132095e+17, 1.288744259172721e+17, 1.288744259213345e+17, 1.288744259252408e+17, 1.288744259293032e+17, 1.288744259332096e+17, 1.288744259372719e+17, 1.288744259413344e+17, 1.288744259452408e+17, 1.288744259493032e+17, 1.288744259532095e+17, 1.288744259572719e+17, 1.288744259613345e+17, 1.288744259652407e+17, 1.288744259693033e+17, 1.288744259732096e+17, 1.288744259772719e+17, 1.288744259813345e+17, 1.288744259852407e+17, 1.288744259893032e+17, 1.288744259932095e+17, 1.288744259972719e+17, 1.288744260013345e+17, 1.288744260052407e+17, 1.288744260093033e+17, 1.288744260132095e+17, 1.288744260172719e+17, 1.288744260213345e+17, 1.288744260252407e+17, 1.288744260293033e+17, 1.288744260332095e+17, 1.288744260372719e+17, 1.288744260413345e+17, 1.288744260452407e+17, 1.288744260493033e+17, 1.288744260532095e+17, 1.288744260572721e+17, 1.288744260613345e+17, 1.288744260652407e+17, 1.288744260693033e+17, 1.288744260732095e+17, 1.288744260772719e+17, 1.288744260813345e+17, 1.288744260852407e+17, 1.288744260893033e+17, 1.288744260932095e+17, 1.288744260972721e+17, 1.288744261013345e+17, 1.288744261052408e+17, 1.288744261093033e+17, 1.288744261132095e+17, 1.288744261172721e+17, 1.288744261213344e+17, 1.288744261252407e+17, 1.288744261293033e+17, 1.288744261332095e+17, 1.288744261372721e+17, 1.288744261413345e+17, 1.288744261452408e+17, 1.288744261493032e+17, 1.288744261532095e+17, 1.288744261572721e+17, 1.288744261613344e+17, 1.288744261652408e+17, 1.288744261693032e+17, 1.288744261732095e+17, 1.288744261772719e+17, 1.288744261813345e+17, 1.288744261852408e+17, 1.288744261893032e+17, 1.288744261932096e+17, 1.288744261972719e+17, 1.288744262013345e+17, 1.288744262052407e+17, 1.288744262093032e+17, 1.288744262132095e+17, 1.288744262172719e+17, 1.288744262213345e+17, 1.288744262252407e+17, 1.288744262293033e+17, 1.288744262332095e+17, 1.288744262372719e+17, 1.288744262413345e+17, 1.288744262452407e+17, 1.288744262493032e+17, 1.288744262532095e+17, 1.288744262572719e+17, 1.288744262613345e+17, 1.288744262652407e+17, 1.288744262693033e+17, 1.288744262732095e+17, 1.288744262772719e+17, 1.288744262813345e+17, 1.288744262852407e+17, 1.288744262893033e+17, 1.288744262932095e+17, 1.288744262972719e+17, 1.288744263013345e+17, 1.288744263052407e+17, 1.288744263093033e+17, 1.288744263132095e+17, 1.288744263172721e+17, 1.288744263213345e+17, 1.288744263252407e+17, 1.288744263293033e+17, 1.288744263332095e+17, 1.288744263372719e+17, 1.288744263413345e+17, 1.288744263452407e+17, 1.288744263493033e+17, 1.288744263532095e+17, 1.288744263572721e+17, 1.288744263613345e+17, 1.288744263652408e+17, 1.288744263693033e+17, 1.288744263732095e+17, 1.288744263772721e+17, 1.288744263813344e+17, 1.288744263852407e+17, 1.288744263893033e+17, 1.288744263932095e+17, 1.288744263972721e+17, 1.288744264013345e+17, 1.288744264052408e+17, 1.288744264093032e+17, 1.288744264132095e+17, 1.288744264172721e+17, 1.288744264213344e+17, 1.288744264252408e+17, 1.288744264293032e+17, 1.288744264332095e+17, 1.288744264372719e+17, 1.288744264413345e+17, 1.288744264452408e+17, 1.288744264493032e+17, 1.288744264532096e+17, 1.288744264572719e+17, 1.288744264613345e+17, 1.288744264652407e+17, 1.288744264693032e+17, 1.288744264732095e+17, 1.288744264772719e+17, 1.288744264813345e+17, 1.288744264852407e+17, 1.288744264893033e+17, 1.288744264932095e+17, 1.288744264972719e+17, 1.288744265013345e+17, 1.288744265052407e+17, 1.288744265093032e+17, 1.288744265132095e+17, 1.288744265172719e+17, 1.288744265213345e+17, 1.288744265252407e+17, 1.288744265293033e+17, 1.288744265332095e+17, 1.288744265372719e+17, 1.288744265413345e+17, 1.288744265452407e+17, 1.288744265493033e+17, 1.288744265532095e+17, 1.288744265572719e+17, 1.288744265613345e+17, 1.288744265652407e+17, 1.288744265693033e+17, 1.288744265732095e+17, 1.288744265772721e+17, 1.288744265813345e+17, 1.288744265852407e+17, 1.288744265893033e+17, 1.288744265932095e+17, 1.288744265972719e+17, 1.288744266013345e+17, 1.288744266052407e+17, 1.288744266093033e+17, 1.288744266132095e+17, 1.288744266172721e+17, 1.288744266213345e+17, 1.288744266252408e+17, 1.288744266293033e+17, 1.288744266332095e+17, 1.288744266372721e+17, 1.288744266413344e+17, 1.288744266452407e+17, 1.288744266493033e+17, 1.288744266532095e+17, 1.288744266572721e+17, 1.288744266613345e+17, 1.288744266652408e+17, 1.288744266693032e+17, 1.288744266732095e+17, 1.288744266772721e+17, 1.288744266813344e+17, 1.288744266852408e+17, 1.288744266893032e+17, 1.288744266932095e+17, 1.288744266972719e+17, 1.288744267013345e+17, 1.288744267052408e+17, 1.288744267093032e+17, 1.288744267132096e+17, 1.288744267172719e+17, 1.288744267213345e+17, 1.288744267252407e+17, 1.288744267293032e+17, 1.288744267332095e+17, 1.288744267372719e+17, 1.288744267413345e+17, 1.288744267452407e+17, 1.288744267493033e+17, 1.288744267532095e+17},
			             {1.288744306213345e+17, 1.288744306252407e+17, 1.288744306293033e+17, 1.288744306332095e+17, 1.288744306372719e+17, 1.288744306413345e+17, 1.288744306452407e+17, 1.288744306493033e+17, 1.288744306532095e+17, 1.288744306572721e+17, 1.288744306613345e+17, 1.288744306652407e+17, 1.288744306693033e+17, 1.288744306732095e+17, 1.288744306772721e+17, 1.288744306813345e+17, 1.288744306852407e+17, 1.288744306893033e+17, 1.288744306932095e+17, 1.288744306972721e+17, 1.288744307013345e+17, 1.288744307052408e+17, 1.288744307093033e+17, 1.288744307132095e+17, 1.288744307172721e+17, 1.288744307213344e+17, 1.288744307252407e+17, 1.288744307293033e+17, 1.288744307332095e+17, 1.288744307372721e+17, 1.288744307413345e+17, 1.288744307452408e+17, 1.288744307493032e+17, 1.288744307532095e+17, 1.288744307572721e+17, 1.288744307613344e+17, 1.288744307652408e+17, 1.288744307693032e+17, 1.288744307732095e+17, 1.288744307772719e+17, 1.288744307813345e+17, 1.288744307852408e+17, 1.288744307893032e+17, 1.288744307932096e+17, 1.288744307972719e+17, 1.288744308013345e+17, 1.288744308052407e+17, 1.288744308093032e+17, 1.288744308132095e+17, 1.288744308172719e+17, 1.288744308213345e+17, 1.288744308252407e+17, 1.288744308293033e+17, 1.288744308332095e+17, 1.288744308372719e+17, 1.288744308413345e+17},
			             {1.288744320652407e+17, 1.288744320693032e+17, 1.288744320732095e+17, 1.288744320772719e+17, 1.288744320813345e+17, 1.288744320852407e+17, 1.288744320893033e+17, 1.288744320932095e+17, 1.288744320972719e+17, 1.288744321013345e+17, 1.288744321052407e+17, 1.288744321093032e+17, 1.288744321132095e+17, 1.288744321172719e+17, 1.288744321213345e+17, 1.288744321252407e+17, 1.288744321293033e+17, 1.288744321332095e+17, 1.288744321372719e+17, 1.288744321413345e+17, 1.288744321452407e+17, 1.288744321493033e+17, 1.288744321532095e+17, 1.288744321572719e+17, 1.288744321613345e+17, 1.288744321652407e+17, 1.288744321693033e+17, 1.288744321732095e+17, 1.288744321772721e+17, 1.288744321813345e+17, 1.288744321852407e+17, 1.288744321893033e+17, 1.288744321932095e+17, 1.288744321972719e+17, 1.288744322013345e+17, 1.288744322052407e+17, 1.288744322093033e+17, 1.288744322132095e+17, 1.288744322172721e+17, 1.288744322213345e+17, 1.288744322252408e+17, 1.288744322293033e+17, 1.288744322332095e+17, 1.288744322372721e+17, 1.288744322413344e+17, 1.288744322452407e+17, 1.288744322493033e+17, 1.288744322532095e+17, 1.288744322572721e+17, 1.288744322613345e+17, 1.288744322652408e+17, 1.288744322693032e+17, 1.288744322732095e+17, 1.288744322772721e+17, 1.288744322813344e+17, 1.288744322852408e+17, 1.288744322893032e+17, 1.288744322932095e+17, 1.288744322972719e+17, 1.288744323013345e+17, 1.288744323052408e+17, 1.288744323093032e+17, 1.288744323132096e+17, 1.288744323172719e+17, 1.288744323213345e+17, 1.288744323252407e+17, 1.288744323293032e+17, 1.288744323332095e+17, 1.288744323372719e+17, 1.288744323413345e+17, 1.288744323452407e+17, 1.288744323493033e+17, 1.288744323532095e+17, 1.288744323572719e+17, 1.288744323613345e+17, 1.288744323652407e+17, 1.288744323693032e+17, 1.288744323732095e+17, 1.288744323772719e+17, 1.288744323813345e+17, 1.288744323852407e+17, 1.288744323893033e+17, 1.288744323932095e+17, 1.288744323972721e+17, 1.288744324013345e+17, 1.288744324052407e+17, 1.288744324093033e+17, 1.288744324132095e+17},
			             {1.288744231693032e+17, 1.288744231732095e+17, 1.288744231772719e+17, 1.288744231813345e+17, 1.288744231852407e+17, 1.288744231893033e+17, 1.288744231932095e+17},
			             {1.288744233813344e+17, 1.288744233852408e+17, 1.288744233893032e+17, 1.288744233932095e+17, 1.288744233972719e+17, 1.288744234013345e+17, 1.288744234052407e+17, 1.288744234093033e+17, 1.288744234132096e+17, 1.288744234172719e+17};
			mask_depths = {{63.1, 64.4}, {63.1, 64.4}, {63.1, 64.4}, {63.1, 64.4}, {63.1, 64.4}, {63.1, 64.4}, {63.1, 64.4}}, {{14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}, {14.0, 26.9}}, {{13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}, {13.9, 23.9}}, {{61.2, 65.0}, {61.2, 65.0}, {61.2, 65.0}, {61.2, 65.0}, {61.2, 65.0}, {61.2, 65.0}, {61.2, 65.0}}, {{55.5, 61.4}, {55.5, 61.4}, {55.5, 61.4}, {55.5, 61.4}, {55.5, 61.4}, {55.5, 61.4}, {55.5, 61.4}}, {{60.3, 62.3}, {60.3, 62.3}, {60.3, 62.3}, {60.3, 62.3}, {60.3, 62.3}}, {{62.7, 65.7}, {62.7, 65.7}, {62.7, 65.7}, {62.7, 65.7}, {62.7, 65.7}, {62.7, 65.7}, {62.7, 65.7}, {62.7, 65.7}}, {{64.2, 65.8}, {64.2, 65.8}, {64.2, 65.8}, {64.2, 65.8}, {64.2, 65.8}, {64.2, 65.8}, {64.2, 65.8}}, {{65.3, 66.6}, {65.3, 66.6}, {65.3, 66.6}, {65.3, 66.6}, {65.3, 66.6}, {65.3, 66.7}, {65.3, 66.7}}, {{64.1, 65.8}, {64.1, 65.8}, {64.1, 65.8}, {64.1, 65.8}, {64.1, 65.8}}, {{68.2, 69.1}, {68.2, 69.2}, {68.2, 69.2}, {68.2, 69.2}, {68.2, 69.2}, {68.2, 69.1}}, {{32.7, 35.8}, {32.7, 35.8}, {32.7, 35.8}, {32.7, 35.8}, {32.7, 35.8}, {32.7, 35.8}}, {{31.9, 34.0}, {31.9, 34.0}, {31.9, 34.0}, {31.9, 34.0}, {31.9, 34.0}}, {{68.1, 72.0}, {67.7, 68.1, 72.1, 72.3}, {67.5, 67.7, 72.2, 72.2}, {67.5, 67.5, 72.3}, {65.4, 67.5, 72.3}, {65.4, 65.4, 72.3}, {65.3, 65.4, 72.3}, {65.3, 72.3}, {65.4, 72.3}, {65.5, 66.1, 72.3}, {66.2, 66.3, 72.3}, {66.4, 72.3}, {66.5, 66.9, 72.2, 72.3}, {67.0, 67.5, 72.2}, {67.6, 67.8, 72.2}, {68.0, 69.2, 72.2}, {69.4, 72.2}}, {{55.4, 58.8}, {53.7, 55.2, 58.8, 59.7}, {53.2, 53.6, 59.9, 60.8}, {53.1, 60.9}, {53.0, 53.1, 61.0, 61.3}, {53.0, 61.3, 61.5}, {52.7, 52.8, 61.6, 61.7}, {52.6, 52.6, 61.7}, {52.3, 52.5, 61.7}, {52.3, 61.7}, {52.3, 61.7}, {52.3, 61.7}, {52.3, 61.7}, {52.3, 61.7}, {52.3, 61.7}, {52.3, 61.7}, {52.3, 61.7}, {52.3, 52.5, 61.7}, {52.6, 52.8, 61.7}, {52.8, 53.1, 61.1, 61.7}, {53.2, 53.8, 60.5, 60.9}, {54.0, 54.4, 59.8, 60.4}, {54.7, 59.8}}, {{53.9, 63.0, 63.9, 65.9}, {53.9, 63.0, 63.8, 66.0}, {53.9, 63.0, 63.8, 66.1}, {53.9, 63.0, 63.7, 66.2, 66.3}, {53.9, 66.5, 66.5}, {53.9, 66.6}, {53.9, 66.6}, {53.9, 66.7}, {53.9, 66.7}, {53.9, 66.6}, {53.9, 66.6}, {53.9, 66.6, 66.6}, {53.9, 66.6}, {53.9, 66.3, 66.4}, {53.9, 66.1}, {53.9, 54.2, 65.5, 65.9}, {54.6, 65.4}, {54.6, 65.3, 65.3}, {54.7, 65.1}, {54.9, 64.8, 65.0}, {54.9, 64.8}, {55.0, 64.7}, {55.0, 64.6}, {55.0, 64.6}, {55.0, 64.5}, {55.0, 64.3}, {55.0, 64.3}, {55.1, 64.3}, {55.1, 64.2, 64.3}, {54.9, 64.2}, {54.9, 64.2}, {54.9, 64.2}, {54.9, 64.2, 64.2}, {54.9, 64.1}, {54.9, 63.9}, {54.9, 63.8}, {54.9, 63.4, 63.7}, {55.0, 55.0, 63.3}, {55.1, 63.1}, {55.2, 63.0}, {55.3, 55.4, 62.7}, {55.8, 62.0}, {56.0, 61.9}, {56.6, 61.9}, {56.7, 61.6}, {56.8, 61.4}, {57.1, 61.1}}, {{54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}, {54.1, 58.6}}, {{62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}, {62.8, 68.4}}, {{52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}, {52.5, 60.6}}, {{52.9, 54.0}, {52.9, 54.0}, {52.9, 54.0}, {52.9, 54.0}, {52.9, 54.0}}, {{56.9, 60.3}, {56.9, 60.3}, {56.9, 60.3}, {56.9, 60.3}, {56.9, 60.3}, {56.9, 60.3}}, {{54.7, 57.8}, {54.7, 57.8}, {54.7, 57.8}, {54.7, 57.8}, {54.7, 57.8}, {54.7, 57.8}, {54.7, 57.8}, {54.7, 57.8}, {54.7, 57.8}}, {{51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}, {51.0, 62.4}}, {{55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}, {55.3, 64.7}}, {{57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}, {57.4, 62.2}}, {{49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}, {49.6, 57.2}}, {{58.5, 64.1}, {58.5, 64.1}, {58.5, 64.1}, {58.5, 64.1}, {58.5, 64.1}, {58.5, 64.1}, {58.5, 64.1}, {58.5, 64.1}, {58.5, 64.1}}, {{55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}, {55.5, 61.8}}, {{60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}, {60.5, 67.8}}, {{68.6, 69.7}, {68.6, 69.7}, {68.6, 69.6}, {68.6, 69.6}, {68.6, 69.6}, {68.6, 69.6}, {68.6, 69.6}, {68.6, 69.6}}, {{68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.7}, {68.0, 69.6}}, {{60.4, 63.1}, {60.4, 63.1}, {60.4, 63.1}, {60.4, 63.1}, {60.4, 63.1}, {60.4, 63.1}, {60.4, 63.1}, {60.4, 63.1}, {60.4, 63.1}, {60.4, 63.1}}, {{64.8, 67.3}, {64.8, 67.3}, {64.8, 67.3}, {64.8, 67.3}, {64.8, 67.3}, {64.8, 67.3}, {64.8, 67.3}, {64.8, 67.3}, {64.8, 67.2}, {64.8, 67.1}}, {{61.4, 63.9}, {61.4, 63.9}, {61.4, 63.9}, {61.4, 63.9}, {61.4, 63.9}, {61.4, 63.9}, {61.4, 63.9}, {61.4, 63.9}, {61.4, 63.9}, {61.4, 63.9}}, {{62.3, 64.9}, {62.3, 64.9}, {62.3, 64.9}, {62.3, 64.9}, {62.3, 64.9}, {62.3, 64.9}, {62.3, 64.9}, {62.3, 64.9}}, {{11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}, {11.2, 31.3}}, {{15.9, 19.7}, {15.6, 20.5}, {14.8, 15.1, 21.2, 21.8}, {14.1, 14.6, 23.0, 25.4}, {13.9, 26.5, 27.0}, {13.4, 27.2}, {13.0, 27.4}, {12.5, 27.6}, {12.4, 12.5, 28.1}, {12.5, 28.3}, {12.2, 28.6}, {12.2, 28.7}, {12.1, 28.8}, {12.0, 28.9}, {11.9, 11.9, 29.0}, {11.8, 29.1}, {11.8, 29.2}, {11.7, 29.4}, {11.6, 29.5}, {11.6, 29.6}, {11.5, 29.6}, {11.5, 29.7}, {11.4, 29.7}, {11.4, 29.7}, {11.4, 29.7}, {11.4, 29.7}, {11.4, 29.7}, {11.3, 29.7}, {11.3, 29.7}, {11.2, 29.3, 29.7}, {11.2, 29.1, 29.2}, {11.2, 29.1}, {11.2, 29.0}, {11.1, 28.9}, {11.1, 28.8}, {11.0, 28.7}, {11.0, 28.6}, {11.0, 28.6}, {11.0, 28.5}, {11.0, 28.4, 28.4}, {11.0, 28.2}, {11.0, 27.6, 28.0}, {11.0, 27.3}, {11.0, 27.1}, {11.0, 26.8}, {11.0, 26.6}, {11.0, 26.4}, {10.9, 11.0, 26.2}, {10.9, 26.1}, {10.9, 25.9}, {10.9, 25.8}, {10.9, 25.7}, {10.9, 25.5}, {10.9, 25.5}, {10.9, 25.4}, {10.9, 25.3}, {10.9, 25.3}, {10.9, 25.2}, {10.9, 25.1, 25.1}, {10.9, 25.1}, {10.9, 25.1}, {10.9, 25.1}, {10.9, 25.1}, {11.0, 25.1}, {11.0, 25.1}, {11.0, 25.1}, {11.1, 25.1}, {11.2, 25.0}, {11.3, 25.0}, {11.3, 25.0}, {11.4, 25.0}, {11.4, 25.0}, {11.5, 25.0}, {11.5, 25.0}, {11.6, 25.0}, {11.7, 25.0}, {11.8, 25.0}, {12.0, 25.0}, {12.1, 25.0}, {12.1, 25.0}, {12.2, 25.0}, {12.3, 25.0}, {12.3, 25.0}, {12.4, 25.0}, {12.4, 25.0}, {12.4, 24.9}, {12.4, 24.9}, {12.4, 24.9}, {12.3, 24.9}, {12.3, 24.9}, {12.2, 24.9}, {12.2, 24.9}, {12.1, 24.9}, {12.1, 24.9}, {12.0, 24.9}, {11.9, 24.9}, {11.9, 24.9}, {11.8, 24.9}, {11.7, 11.8, 24.9}, {11.7, 24.9}, {11.7, 24.9}, {11.9, 24.9}, {11.8, 24.9}, {11.7, 24.9}, {11.6, 24.9}, {11.6, 24.9}, {11.5, 24.9}, {11.4, 24.9}, {11.3, 24.9}, {11.2, 24.9}, {11.2, 24.9}, {11.1, 24.9}, {11.1, 24.9}, {11.1, 24.9}, {11.0, 24.9}, {11.0, 24.9}, {11.0, 24.9}, {11.0, 24.9}, {11.0, 24.9}, {11.0, 24.9}, {11.0, 24.9}, {11.0, 24.9, 25.0}, {11.0, 25.0}, {11.0, 25.0}, {11.0, 25.0}, {11.0, 25.0}, {11.0, 25.0}, {11.0, 25.0}, {11.0, 25.0}, {11.0, 11.1, 25.0}, {11.1, 25.1}, {11.1, 25.1}, {11.1, 25.1}, {11.2, 25.1}, {11.2, 25.1}, {11.3, 25.1}, {11.3, 25.1}, {11.4, 25.1}, {11.4, 25.1}, {11.5, 25.1}, {11.6, 25.1}, {11.8, 25.2}, {11.9, 25.2}, {11.9, 25.2}, {12.0, 25.2}, {12.2, 25.2}, {12.4, 25.3}, {12.5, 25.3}, {12.6, 25.3}, {12.7, 25.3}, {12.8, 25.3}, {12.9, 25.4}, {13.0, 25.4}, {13.1, 25.4}, {13.2, 25.4}, {13.3, 25.4}, {13.3, 25.5}, {13.4, 25.5}, {13.5, 25.5}, {13.5, 25.5}, {13.6, 25.6}, {13.7, 25.6}, {13.7, 25.6}, {13.8, 25.6}, {13.8, 25.6}, {13.8, 25.6}, {13.8, 25.5}, {13.8, 25.5}, {13.9, 25.5}, {13.8, 25.5}, {13.8, 25.5}, {13.7, 25.5}, {13.7, 25.5}, {13.7, 25.5}, {13.6, 25.5}, {13.6, 25.5}, {13.5, 25.5}, {13.4, 25.5}, {13.3, 25.5}, {13.3, 25.5}, {13.2, 25.5}, {13.1, 25.5}, {12.9, 25.5}, {12.8, 25.5}, {12.8, 25.5}, {12.7, 25.5}, {12.6, 25.5}, {12.6, 25.5}, {12.5, 25.5}, {12.5, 25.6}, {12.4, 25.6}, {12.4, 25.6}, {12.3, 25.6}, {12.3, 25.7}, {12.2, 25.7}, {12.2, 25.8}, {12.1, 25.8}, {12.1, 25.9}, {12.0, 25.9}, {11.9, 12.0, 26.1}, {11.8, 26.2}, {11.8, 26.4}, {11.7, 26.5}, {11.6, 26.7}, {11.6, 26.8}, {11.6, 27.0}, {11.6, 27.1}, {11.6, 27.3}, {11.5, 27.7}, {11.5, 28.1}, {11.5, 28.4}, {11.5, 28.7, 29.1}, {11.5, 29.4}, {11.5, 29.6}, {11.5, 29.7}, {11.5, 29.9}, {11.6, 30.1}, {11.6, 30.3}, {11.6, 30.5}, {11.7, 30.7}, {11.7, 30.8, 31.0}, {11.8, 31.1}, {11.8, 31.2}, {11.9, 31.4}, {12.0, 31.5, 31.8}, {12.0, 31.8}, {12.1, 31.8}, {12.1, 31.8}, {12.2, 31.8}, {12.2, 31.7}, {12.2, 31.7}, {12.3, 31.7}, {12.3, 31.7}, {12.3, 31.7}, {12.4, 31.7}, {12.5, 31.7}, {12.6, 31.6}, {12.7, 31.6}, {12.8, 31.6}, {12.9, 31.6}, {13.0, 31.6}, {13.1, 31.6}, {13.3, 31.6}, {13.4, 31.6}, {13.5, 31.6}, {13.7, 31.6}, {13.8, 31.5}, {14.0, 31.5}, {14.1, 31.0}, {14.2, 31.1}, {14.4, 31.1}, {14.5, 31.1}, {14.6, 30.9}, {14.7, 30.6}, {15.0, 30.2}, {15.2, 29.9}, {15.5, 29.6}, {15.8, 29.2}, {15.9, 28.9}, {16.1, 16.4, 28.1}, {16.6, 27.4}, {16.8, 26.7}, {17.1, 26.2}, {17.5, 25.1}, {18.1, 24.0}, {18.7, 22.9}}, {{9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}, {9.8, 31.9}}, {{11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}, {11.6, 34.4}}, {{61.2, 63.2}, {61.2, 63.2}, {61.2, 63.2}, {61.2, 63.2}, {61.2, 63.2}, {61.2, 63.2}, {61.2, 63.2}}, {{64.2, 65.7}, {64.2, 65.7}, {64.2, 65.7}, {64.2, 65.7}, {64.2, 65.7}, {64.2, 65.7}, {64.2, 65.7}, {64.2, 65.7}, {64.2, 65.7}, {64.2, 65.7}};
		}
	}
}
