netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 27;
			channels = 4;
			categories = 108;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  13.0, 39.8, 39.9, 39.2, 39.1, 36.9, 38.9, 39.9, 40.2, 38.4, 37.6, 37.4, 37.4, 37.4, 37.5, 36.3, 36.4, 37.2, 37.0, 37.6, 36.5, 36.8, 30.0, 35.9, 21.9, 41.8, 42.3;
			max_depth =  55.4, 42.9, 41.6, 41.0, 40.4, 40.2, 40.0, 40.9, 41.0, 39.6, 38.7, 38.5, 38.5, 38.5, 38.5, 37.7, 38.1, 38.0, 38.0, 38.6, 38.3, 38.8, 36.1, 38.8, 31.8, 44.9, 45.6;
			start_time = 129799100817695744, 129799100934102016, 129799101572695808, 129799101677070720, 129799101701133184, 129799101765352064, 129799101797539456, 129799101825664512, 129799101837695744, 129799101966289536, 129799101978320768, 129799102150977024, 129799102175039488, 129799102215195776, 129799102243320832, 129799102476289536, 129799102492383232, 129799102516445696, 129799102536445696, 129799102596758272, 129799102693164416, 129799102809570816, 129799102905976960, 129799102938164480, 129799117242851968, 129799106066445824, 129799106295352064;
			end_time = 129799118664570752, 129799100970195712, 129799101588789504, 129799101697070720, 129799101713164544, 129799101789570816, 129799101805664512, 129799101833633152, 129799101845820672, 129799101974258304, 129799101990352000, 129799102158945792, 129799102179102080, 129799102223320832, 129799102247383168, 129799102484258176, 129799102512383232, 129799102528476928, 129799102548477056, 129799102608789504, 129799102713164544, 129799102845664512, 129799102922070784, 129799102950195712, 129799117295195776, 129799106094570752, 129799106335664512;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27;
			region_name = "Layer1","Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21","Layer22","Layer23","Layer24","Layer25","Layer26";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "0", "0", "0", "0", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "200", "333";
			region_channels = 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15;
			mask_times = {1.297991008176957e+17, 1.297991008216019e+17, 1.297991008256645e+17, 1.29799100829727e+17, 1.297991008337894e+17, 1.297991008376957e+17, 1.297991008417583e+17, 1.297991008458207e+17, 1.297991008497271e+17, 1.297991008537894e+17, 1.29799100857852e+17, 1.297991008619145e+17, 1.297991008658207e+17, 1.297991008698833e+17, 1.297991008739457e+17, 1.29799100877852e+17, 1.297991008819146e+17, 1.29799100885977e+17, 1.297991008898833e+17, 1.297991008939457e+17, 1.297991008980082e+17, 1.297991009020708e+17, 1.29799100905977e+17, 1.297991009100396e+17, 1.29799100914102e+17, 1.297991009180083e+17, 1.297991009220708e+17, 1.297991009261332e+17, 1.297991009300396e+17, 1.29799100934102e+17, 1.297991009381645e+17, 1.297991009420708e+17, 1.297991009461332e+17, 1.297991009501957e+17, 1.297991009542583e+17, 1.297991009581645e+17, 1.297991009622269e+17, 1.297991009662895e+17, 1.297991009701957e+17, 1.297991009742583e+17, 1.297991009783208e+17, 1.297991009823832e+17, 1.297991009862895e+17, 1.29799100990352e+17, 1.297991009944145e+17, 1.297991009983206e+17, 1.297991010023832e+17, 1.297991010064458e+17, 1.29799101010352e+17, 1.297991010144146e+17, 1.297991010184769e+17, 1.297991010225395e+17, 1.297991010264458e+17, 1.297991010305082e+17, 1.297991010345708e+17, 1.297991010384769e+17, 1.297991010425395e+17, 1.297991010466021e+17, 1.297991010506644e+17, 1.297991010545708e+17, 1.297991010586332e+17, 1.297991010626957e+17, 1.29799101066602e+17, 1.297991010706644e+17, 1.29799101074727e+17, 1.297991010786332e+17, 1.297991010826958e+17, 1.297991010867583e+17, 1.297991010908207e+17, 1.29799101094727e+17, 1.297991010987895e+17, 1.29799101102852e+17, 1.297991011067583e+17, 1.297991011108207e+17, 1.297991011148832e+17, 1.297991011187895e+17, 1.29799101122852e+17, 1.297991011269144e+17, 1.297991011308207e+17, 1.297991011348832e+17, 1.297991011389458e+17, 1.297991011430083e+17, 1.297991011469146e+17, 1.29799101150977e+17, 1.297991011550395e+17, 1.297991011589458e+17, 1.297991011630081e+17, 1.297991011670707e+17, 1.297991011711333e+17, 1.297991011750395e+17, 1.297991011791021e+17, 1.297991011831645e+17, 1.297991011870707e+17, 1.297991011911333e+17, 1.297991011951956e+17, 1.29799101199102e+17, 1.297991012031645e+17, 1.29799101207227e+17, 1.297991012112896e+17, 1.297991012151958e+17, 1.297991012192582e+17, 1.297991012233208e+17, 1.29799101227227e+17, 1.297991012312895e+17, 1.297991012353519e+17, 1.297991012394145e+17, 1.297991012433208e+17, 1.297991012473833e+17, 1.297991012514458e+17, 1.297991012553519e+17, 1.297991012594145e+17, 1.29799101263477e+17, 1.297991012673832e+17, 1.297991012714458e+17, 1.297991012755082e+17, 1.297991012795707e+17, 1.297991012834771e+17, 1.297991012875395e+17, 1.297991012916019e+17, 1.297991012955082e+17, 1.297991012995707e+17, 1.297991013036333e+17, 1.297991013075395e+17, 1.29799101311602e+17, 1.297991013156645e+17, 1.297991013195708e+17, 1.297991013236333e+17, 1.297991013276957e+17, 1.297991013317582e+17, 1.297991013356645e+17, 1.29799101339727e+17, 1.297991013437896e+17, 1.297991013476957e+17, 1.297991013517582e+17, 1.297991013558208e+17, 1.297991013598833e+17, 1.297991013637894e+17, 1.29799101367852e+17, 1.297991013719145e+17, 1.297991013758208e+17, 1.297991013798833e+17, 1.297991013839457e+17, 1.29799101387852e+17, 1.297991013919145e+17, 1.29799101395977e+17, 1.297991014000396e+17, 1.297991014039457e+17, 1.297991014080083e+17, 1.297991014120708e+17, 1.297991014159771e+17, 1.297991014200394e+17, 1.29799101424102e+17, 1.297991014281645e+17, 1.297991014320707e+17, 1.297991014361332e+17, 1.297991014401958e+17, 1.29799101444102e+17, 1.297991014481646e+17, 1.297991014522269e+17, 1.297991014561332e+17, 1.297991014601958e+17, 1.297991014642582e+17, 1.297991014683208e+17, 1.297991014722269e+17, 1.297991014762895e+17, 1.29799101480352e+17, 1.297991014842583e+17, 1.297991014883208e+17, 1.297991014923832e+17, 1.297991014962895e+17, 1.29799101500352e+17, 1.297991015044145e+17, 1.297991015083208e+17, 1.297991015123832e+17, 1.297991015164457e+17, 1.297991015205083e+17, 1.297991015244145e+17, 1.297991015284769e+17, 1.297991015325395e+17, 1.297991015364457e+17, 1.297991015405083e+17, 1.297991015445708e+17, 1.297991015486332e+17, 1.297991015525395e+17, 1.29799101556602e+17, 1.297991015606644e+17, 1.297991015645708e+17, 1.297991015686332e+17, 1.297991015726958e+17, 1.29799101576602e+17, 1.297991015806646e+17, 1.29799101584727e+17, 1.297991015887895e+17, 1.297991015926958e+17, 1.297991015967581e+17, 1.297991016008207e+17, 1.29799101604727e+17, 1.297991016087895e+17, 1.297991016128521e+17, 1.297991016169146e+17, 1.297991016208207e+17, 1.297991016248833e+17, 1.297991016289457e+17, 1.29799101632852e+17, 1.297991016369144e+17, 1.29799101640977e+17, 1.297991016448833e+17, 1.297991016489458e+17, 1.297991016530083e+17, 1.297991016570707e+17, 1.29799101660977e+17, 1.297991016650395e+17, 1.29799101669102e+17, 1.297991016730083e+17, 1.297991016770707e+17, 1.297991016811332e+17, 1.297991016850396e+17, 1.29799101689102e+17, 1.297991016931645e+17, 1.297991016970707e+17, 1.297991017011332e+17, 1.297991017051958e+17, 1.297991017092582e+17, 1.297991017131645e+17, 1.29799101717227e+17, 1.297991017212895e+17, 1.297991017251958e+17, 1.297991017292582e+17, 1.297991017333207e+17, 1.297991017373833e+17, 1.297991017412895e+17, 1.297991017453521e+17, 1.297991017494145e+17, 1.297991017533207e+17, 1.297991017573833e+17, 1.297991017614458e+17, 1.297991017653521e+17, 1.297991017694145e+17, 1.29799101773477e+17, 1.297991017775396e+17, 1.297991017814458e+17, 1.297991017855082e+17, 1.297991017895708e+17, 1.29799101793477e+17, 1.297991017975395e+17, 1.29799101801602e+17, 1.297991018056645e+17, 1.297991018095708e+17, 1.297991018136333e+17, 1.297991018176957e+17, 1.297991018216019e+17, 1.297991018256645e+17, 1.29799101829727e+17, 1.297991018336332e+17, 1.297991018376957e+17, 1.297991018417583e+17, 1.297991018458207e+17, 1.297991018497271e+17, 1.297991018537894e+17, 1.29799101857852e+17, 1.297991018617583e+17, 1.297991018658207e+17, 1.297991018698833e+17, 1.297991018737894e+17, 1.29799101877852e+17, 1.297991018819145e+17, 1.297991018858208e+17, 1.297991018898833e+17, 1.297991018939457e+17, 1.297991018980082e+17, 1.297991019019145e+17, 1.29799101905977e+17, 1.297991019100396e+17, 1.297991019139457e+17, 1.297991019180082e+17, 1.297991019220708e+17, 1.297991019261332e+17, 1.297991019300396e+17, 1.29799101934102e+17, 1.297991019381645e+17, 1.297991019420708e+17, 1.297991019461332e+17, 1.297991019501957e+17, 1.29799101954102e+17, 1.297991019581645e+17, 1.297991019622269e+17, 1.297991019662895e+17, 1.297991019701957e+17, 1.297991019742583e+17, 1.297991019783208e+17, 1.297991019822271e+17, 1.297991019862895e+17, 1.29799101990352e+17, 1.297991019944145e+17, 1.297991019983206e+17, 1.297991020023832e+17, 1.297991020064458e+17, 1.29799102010352e+17, 1.297991020144146e+17, 1.297991020184771e+17, 1.297991020223832e+17, 1.297991020264458e+17, 1.297991020305082e+17, 1.297991020345708e+17, 1.297991020384769e+17, 1.297991020425395e+17, 1.29799102046602e+17, 1.297991020505083e+17, 1.297991020545708e+17, 1.297991020586333e+17, 1.297991020625395e+17, 1.29799102066602e+17, 1.297991020706644e+17, 1.297991020745708e+17, 1.297991020786332e+17, 1.297991020826957e+17, 1.297991020867583e+17, 1.297991020906644e+17, 1.29799102094727e+17, 1.297991020987895e+17, 1.297991021026957e+17, 1.297991021067583e+17, 1.297991021108207e+17, 1.297991021148832e+17, 1.297991021187895e+17, 1.29799102122852e+17, 1.297991021269144e+17, 1.297991021308207e+17, 1.297991021348832e+17, 1.297991021389458e+17, 1.29799102142852e+17, 1.297991021469146e+17, 1.29799102150977e+17, 1.297991021550395e+17, 1.297991021589458e+17, 1.297991021630083e+17, 1.297991021670707e+17, 1.29799102170977e+17, 1.297991021750395e+17, 1.297991021791021e+17, 1.297991021831645e+17, 1.297991021870707e+17, 1.297991021911333e+17, 1.297991021951958e+17, 1.29799102199102e+17, 1.297991022031645e+17, 1.29799102207227e+17, 1.297991022111333e+17, 1.297991022151958e+17, 1.297991022192582e+17, 1.297991022233208e+17, 1.29799102227227e+17, 1.297991022312895e+17, 1.297991022353521e+17, 1.297991022392582e+17, 1.297991022433208e+17, 1.297991022473832e+17, 1.297991022512896e+17, 1.297991022553519e+17, 1.297991022594145e+17, 1.297991022633208e+17, 1.297991022673832e+17, 1.297991022714458e+17, 1.297991022755084e+17, 1.297991022794145e+17, 1.29799102283477e+17, 1.297991022875395e+17, 1.297991022914458e+17, 1.297991022955082e+17, 1.297991022995707e+17, 1.297991023036333e+17, 1.297991023075395e+17, 1.29799102311602e+17, 1.297991023156645e+17, 1.297991023195707e+17, 1.297991023236333e+17, 1.297991023276957e+17, 1.29799102331602e+17, 1.297991023356645e+17, 1.29799102339727e+17, 1.297991023437896e+17, 1.297991023476957e+17, 1.297991023517582e+17, 1.297991023558208e+17, 1.29799102359727e+17, 1.297991023637894e+17, 1.29799102367852e+17, 1.297991023719145e+17, 1.297991023758208e+17, 1.297991023798833e+17, 1.297991023839457e+17, 1.29799102387852e+17, 1.297991023919145e+17, 1.29799102395977e+17, 1.297991023998831e+17, 1.297991024039457e+17, 1.297991024080083e+17, 1.297991024120707e+17, 1.297991024159771e+17, 1.297991024200396e+17, 1.29799102424102e+17, 1.297991024280083e+17, 1.297991024320707e+17, 1.297991024361332e+17, 1.297991024400394e+17, 1.29799102444102e+17, 1.297991024481645e+17, 1.297991024520708e+17, 1.297991024561332e+17, 1.297991024601958e+17, 1.297991024642582e+17, 1.297991024681645e+17, 1.297991024722269e+17, 1.297991024762895e+17, 1.297991024801957e+17, 1.297991024842582e+17, 1.297991024883208e+17, 1.297991024923832e+17, 1.297991024962895e+17, 1.29799102500352e+17, 1.297991025044145e+17, 1.297991025083208e+17, 1.297991025123832e+17, 1.297991025164457e+17, 1.29799102520352e+17, 1.297991025244145e+17, 1.297991025284769e+17, 1.297991025325395e+17, 1.297991025364457e+17, 1.297991025405083e+17, 1.297991025445708e+17, 1.297991025484771e+17, 1.297991025525395e+17, 1.29799102556602e+17, 1.297991025606644e+17, 1.297991025645708e+17, 1.297991025686332e+17, 1.297991025726958e+17, 1.29799102576602e+17, 1.297991025806646e+17, 1.29799102584727e+17, 1.297991025886332e+17, 1.297991025926958e+17, 1.297991025967583e+17, 1.297991026008207e+17, 1.29799102604727e+17, 1.297991026087895e+17, 1.29799102612852e+17, 1.297991026167583e+17, 1.297991026208207e+17, 1.297991026248833e+17, 1.297991026287895e+17, 1.29799102632852e+17, 1.297991026369146e+17, 1.297991026408207e+17, 1.297991026448833e+17, 1.297991026489457e+17, 1.297991026530083e+17, 1.297991026569144e+17, 1.29799102660977e+17, 1.297991026650395e+17, 1.297991026689457e+17, 1.297991026730083e+17, 1.297991026770708e+17, 1.297991026811332e+17, 1.297991026850395e+17, 1.29799102689102e+17, 1.297991026931644e+17, 1.297991026970707e+17, 1.297991027011332e+17, 1.297991027051958e+17, 1.29799102709102e+17, 1.297991027131645e+17, 1.29799102717227e+17, 1.297991027212895e+17, 1.297991027251958e+17, 1.297991027292582e+17, 1.297991027333207e+17, 1.29799102737227e+17, 1.297991027412895e+17, 1.297991027453521e+17, 1.297991027494145e+17, 1.297991027533207e+17, 1.297991027573833e+17, 1.297991027614458e+17, 1.297991027653519e+17, 1.297991027694145e+17, 1.29799102773477e+17, 1.297991027773833e+17, 1.297991027814458e+17, 1.297991027855082e+17, 1.297991027895708e+17, 1.29799102793477e+17, 1.297991027975395e+17, 1.29799102801602e+17, 1.297991028055082e+17, 1.297991028095708e+17, 1.297991028136332e+17, 1.297991028175396e+17, 1.29799102821602e+17, 1.297991028256645e+17, 1.297991028295708e+17, 1.297991028336332e+17, 1.297991028376957e+17, 1.297991028417583e+17, 1.297991028456645e+17, 1.29799102849727e+17, 1.297991028537896e+17, 1.297991028576957e+17, 1.297991028617583e+17, 1.297991028658207e+17, 1.297991028698833e+17, 1.297991028737894e+17, 1.29799102877852e+17, 1.297991028819145e+17, 1.297991028858208e+17, 1.297991028898833e+17, 1.297991028939457e+17, 1.29799102897852e+17, 1.297991029019145e+17, 1.29799102905977e+17, 1.297991029100396e+17, 1.297991029139457e+17, 1.297991029180082e+17, 1.297991029220708e+17, 1.29799102925977e+17, 1.297991029300394e+17, 1.29799102934102e+17, 1.297991029381645e+17, 1.297991029420708e+17, 1.297991029461332e+17, 1.297991029501957e+17, 1.29799102954102e+17, 1.297991029581645e+17, 1.297991029622269e+17, 1.297991029661332e+17, 1.297991029701957e+17, 1.297991029742583e+17, 1.297991029783208e+17, 1.297991029822271e+17, 1.297991029862895e+17, 1.29799102990352e+17, 1.297991029942583e+17, 1.297991029983208e+17, 1.297991030023832e+17, 1.297991030062895e+17, 1.29799103010352e+17, 1.297991030144146e+17, 1.297991030183208e+17, 1.297991030223832e+17, 1.297991030264458e+17, 1.297991030305082e+17, 1.297991030344145e+17, 1.297991030384771e+17, 1.297991030425395e+17, 1.297991030464458e+17, 1.297991030505083e+17, 1.297991030545708e+17, 1.297991030586332e+17, 1.297991030625395e+17, 1.29799103066602e+17, 1.297991030706644e+17, 1.297991030745708e+17, 1.297991030786333e+17, 1.297991030826957e+17, 1.297991030866021e+17, 1.297991030906644e+17, 1.297991030947269e+17, 1.297991030987895e+17, 1.297991031026957e+17, 1.297991031067583e+17, 1.297991031108209e+17, 1.29799103114727e+17, 1.297991031187895e+17, 1.29799103122852e+17, 1.297991031269144e+17, 1.297991031308207e+17, 1.297991031348832e+17, 1.297991031389458e+17, 1.29799103142852e+17, 1.297991031469146e+17, 1.29799103150977e+17, 1.297991031548832e+17, 1.297991031589458e+17, 1.297991031630083e+17, 1.297991031670707e+17, 1.29799103170977e+17, 1.297991031750395e+17, 1.297991031791021e+17, 1.297991031830083e+17, 1.297991031870707e+17, 1.297991031911333e+17, 1.297991031950395e+17, 1.29799103199102e+17, 1.297991032031645e+17, 1.297991032070707e+17, 1.297991032111333e+17, 1.297991032151958e+17, 1.297991032192582e+17, 1.297991032231645e+17, 1.29799103227227e+17, 1.297991032312895e+17, 1.297991032351956e+17, 1.297991032392582e+17, 1.297991032433208e+17, 1.297991032473832e+17, 1.297991032512896e+17, 1.297991032553521e+17, 1.297991032594144e+17, 1.297991032633208e+17, 1.297991032673832e+17, 1.297991032714458e+17, 1.297991032753519e+17, 1.297991032794145e+17, 1.29799103283477e+17, 1.297991032875395e+17, 1.297991032914458e+17, 1.297991032955082e+17, 1.297991032995707e+17, 1.29799103303477e+17, 1.297991033075395e+17, 1.29799103311602e+17, 1.297991033156645e+17, 1.297991033195707e+17, 1.297991033236333e+17, 1.297991033276957e+17, 1.297991033316019e+17, 1.297991033356645e+17, 1.29799103339727e+17, 1.297991033436333e+17, 1.297991033476957e+17, 1.297991033517582e+17, 1.297991033558208e+17, 1.29799103359727e+17, 1.297991033637894e+17, 1.29799103367852e+17, 1.297991033717582e+17, 1.297991033758208e+17, 1.297991033798833e+17, 1.297991033837896e+17, 1.29799103387852e+17, 1.297991033919145e+17, 1.297991033958208e+17, 1.297991033998833e+17, 1.297991034039457e+17, 1.297991034080083e+17, 1.297991034119145e+17, 1.297991034159771e+17, 1.297991034200396e+17, 1.297991034239457e+17, 1.297991034280083e+17, 1.297991034320707e+17, 1.297991034361332e+17, 1.297991034400396e+17, 1.29799103444102e+17, 1.297991034481645e+17, 1.297991034520708e+17, 1.297991034561332e+17, 1.297991034601957e+17, 1.29799103464102e+17, 1.297991034681645e+17, 1.297991034722269e+17, 1.297991034762895e+17, 1.297991034801958e+17, 1.297991034842582e+17, 1.297991034883208e+17, 1.297991034922269e+17, 1.297991034962894e+17, 1.29799103500352e+17, 1.297991035044145e+17, 1.297991035083208e+17, 1.297991035123834e+17, 1.297991035164457e+17, 1.29799103520352e+17, 1.297991035244145e+17, 1.297991035284769e+17, 1.297991035323832e+17, 1.297991035364457e+17, 1.297991035405083e+17, 1.297991035445708e+17, 1.297991035484771e+17, 1.297991035525395e+17, 1.29799103556602e+17, 1.297991035605083e+17, 1.297991035645708e+17, 1.297991035686332e+17, 1.297991035725395e+17, 1.29799103576602e+17, 1.297991035806646e+17, 1.297991035845708e+17, 1.297991035886332e+17, 1.297991035926958e+17, 1.297991035967583e+17, 1.297991036006644e+17, 1.29799103604727e+17, 1.297991036087895e+17, 1.297991036126958e+17, 1.297991036167583e+17, 1.297991036208207e+17, 1.297991036248832e+17, 1.297991036287895e+17, 1.29799103632852e+17, 1.297991036369146e+17, 1.297991036408207e+17, 1.297991036448833e+17, 1.297991036489457e+17, 1.297991036528521e+17, 1.297991036569146e+17, 1.297991036609769e+17, 1.297991036650395e+17, 1.297991036689457e+17, 1.297991036730083e+17, 1.297991036770708e+17, 1.29799103680977e+17, 1.297991036850395e+17, 1.29799103689102e+17, 1.297991036931644e+17, 1.297991036970708e+17, 1.297991037011332e+17, 1.297991037051958e+17, 1.29799103709102e+17, 1.297991037131645e+17, 1.29799103717227e+17, 1.297991037211332e+17, 1.297991037251958e+17, 1.297991037292582e+17, 1.297991037333207e+17, 1.29799103737227e+17, 1.297991037412895e+17, 1.297991037453521e+17, 1.297991037492582e+17, 1.297991037533207e+17, 1.297991037573833e+17, 1.297991037612895e+17, 1.297991037653519e+17, 1.297991037694145e+17, 1.297991037733207e+17, 1.297991037773833e+17, 1.297991037814458e+17, 1.297991037855082e+17, 1.297991037894145e+17, 1.29799103793477e+17, 1.297991037975395e+17, 1.297991038014458e+17, 1.297991038055082e+17, 1.297991038095708e+17, 1.297991038136333e+17, 1.297991038175396e+17, 1.29799103821602e+17, 1.297991038256645e+17, 1.297991038295708e+17, 1.297991038336332e+17, 1.297991038376957e+17, 1.29799103841602e+17, 1.297991038456645e+17, 1.29799103849727e+17, 1.297991038537896e+17, 1.297991038576957e+17, 1.297991038617583e+17, 1.297991038658207e+17, 1.29799103869727e+17, 1.297991038737896e+17, 1.29799103877852e+17, 1.297991038819145e+17, 1.297991038858207e+17, 1.297991038898833e+17, 1.297991038939457e+17, 1.29799103897852e+17, 1.297991039019145e+17, 1.29799103905977e+17, 1.297991039098833e+17, 1.297991039139459e+17, 1.297991039180082e+17, 1.297991039220708e+17, 1.29799103925977e+17, 1.297991039300394e+17, 1.29799103934102e+17, 1.297991039380082e+17, 1.297991039420708e+17, 1.297991039461332e+17, 1.297991039500396e+17, 1.29799103954102e+17, 1.297991039581645e+17, 1.297991039620708e+17, 1.297991039661332e+17, 1.297991039701957e+17, 1.297991039742583e+17, 1.297991039781645e+17, 1.297991039822271e+17, 1.297991039862895e+17, 1.297991039901957e+17, 1.297991039942583e+17, 1.297991039983208e+17, 1.297991040023832e+17, 1.297991040062895e+17, 1.29799104010352e+17, 1.297991040144145e+17, 1.297991040183208e+17, 1.297991040223832e+17, 1.297991040264458e+17, 1.29799104030352e+17, 1.297991040344145e+17, 1.297991040384771e+17, 1.297991040425395e+17, 1.297991040464458e+17, 1.297991040505082e+17, 1.297991040545708e+17, 1.297991040584771e+17, 1.297991040625395e+17, 1.29799104066602e+17, 1.297991040706646e+17, 1.297991040745708e+17, 1.297991040786333e+17, 1.297991040826957e+17, 1.29799104086602e+17, 1.297991040906644e+17, 1.297991040947269e+17, 1.297991040986333e+17, 1.297991041026957e+17, 1.297991041067583e+17, 1.297991041108209e+17, 1.29799104114727e+17, 1.297991041187895e+17, 1.29799104122852e+17, 1.297991041267583e+17, 1.297991041308207e+17, 1.297991041348832e+17, 1.297991041387895e+17, 1.29799104142852e+17, 1.297991041469146e+17, 1.297991041508207e+17, 1.297991041548832e+17, 1.297991041589458e+17, 1.297991041630083e+17, 1.297991041669144e+17, 1.29799104170977e+17, 1.297991041750395e+17, 1.297991041789458e+17, 1.297991041830083e+17, 1.297991041870707e+17, 1.297991041911333e+17, 1.297991041950395e+17, 1.29799104199102e+17, 1.297991042031645e+17, 1.297991042070707e+17, 1.297991042111333e+17, 1.297991042151958e+17, 1.297991042191021e+17, 1.297991042231645e+17, 1.29799104227227e+17, 1.297991042312895e+17, 1.297991042351956e+17, 1.297991042392582e+17, 1.297991042433208e+17, 1.29799104247227e+17, 1.297991042512895e+17, 1.297991042553521e+17, 1.297991042594144e+17, 1.297991042633208e+17, 1.297991042673832e+17, 1.297991042714458e+17, 1.297991042753521e+17, 1.297991042794145e+17, 1.29799104283477e+17, 1.297991042873832e+17, 1.297991042914458e+17, 1.297991042955082e+17, 1.297991042995707e+17, 1.29799104303477e+17, 1.297991043075395e+17, 1.29799104311602e+17, 1.297991043155084e+17, 1.297991043195707e+17, 1.297991043236333e+17, 1.297991043275395e+17, 1.297991043316019e+17, 1.297991043356645e+17, 1.297991043395707e+17, 1.297991043436333e+17, 1.297991043476957e+17, 1.297991043517582e+17, 1.297991043556645e+17, 1.29799104359727e+17, 1.297991043637894e+17, 1.297991043676957e+17, 1.297991043717582e+17, 1.297991043758208e+17, 1.297991043798833e+17, 1.297991043837896e+17, 1.29799104387852e+17, 1.297991043919145e+17, 1.297991043958208e+17, 1.297991043998833e+17, 1.297991044039457e+17, 1.29799104407852e+17, 1.297991044119145e+17, 1.29799104415977e+17, 1.297991044200396e+17, 1.297991044239457e+17, 1.297991044280083e+17, 1.297991044320708e+17, 1.29799104435977e+17, 1.297991044400396e+17, 1.29799104444102e+17, 1.297991044481645e+17, 1.297991044520707e+17, 1.297991044561332e+17, 1.297991044601957e+17, 1.29799104464102e+17, 1.297991044681645e+17, 1.297991044722271e+17, 1.297991044761332e+17, 1.297991044801958e+17, 1.297991044842582e+17, 1.297991044883208e+17, 1.297991044922269e+17, 1.297991044962894e+17, 1.29799104500352e+17, 1.297991045042582e+17, 1.297991045083208e+17, 1.297991045123834e+17, 1.297991045162895e+17, 1.29799104520352e+17, 1.297991045244145e+17, 1.297991045283208e+17, 1.297991045323832e+17, 1.297991045364457e+17, 1.297991045405083e+17, 1.297991045444145e+17, 1.297991045484771e+17, 1.297991045525395e+17, 1.297991045564457e+17, 1.297991045605083e+17, 1.297991045645708e+17, 1.297991045686332e+17, 1.297991045725395e+17, 1.29799104576602e+17, 1.297991045806644e+17, 1.297991045845708e+17, 1.297991045886332e+17, 1.297991045926958e+17, 1.29799104596602e+17, 1.297991046006644e+17, 1.29799104604727e+17, 1.297991046087895e+17, 1.297991046126958e+17, 1.297991046167583e+17, 1.297991046208207e+17, 1.29799104624727e+17, 1.297991046287895e+17, 1.29799104632852e+17, 1.297991046369146e+17, 1.297991046408207e+17, 1.297991046448833e+17, 1.297991046489458e+17, 1.29799104652852e+17, 1.297991046569146e+17, 1.297991046609769e+17, 1.297991046648833e+17, 1.297991046689457e+17, 1.297991046730083e+17, 1.297991046770708e+17, 1.29799104680977e+17, 1.297991046850395e+17, 1.297991046891021e+17, 1.297991046930083e+17, 1.297991046970707e+17, 1.297991047011332e+17, 1.297991047050395e+17, 1.29799104709102e+17, 1.297991047131645e+17, 1.297991047170708e+17, 1.297991047211332e+17, 1.297991047251958e+17, 1.297991047292582e+17, 1.297991047331644e+17, 1.29799104737227e+17, 1.297991047412895e+17, 1.297991047451958e+17, 1.297991047492582e+17, 1.297991047533207e+17, 1.297991047573833e+17, 1.297991047612895e+17, 1.297991047653519e+17, 1.297991047694145e+17, 1.297991047733207e+17, 1.297991047773833e+17, 1.297991047814458e+17, 1.297991047853521e+17, 1.297991047894145e+17, 1.29799104793477e+17, 1.297991047975395e+17, 1.297991048014458e+17, 1.297991048055082e+17, 1.297991048095708e+17, 1.29799104813477e+17, 1.297991048175395e+17, 1.29799104821602e+17, 1.297991048256644e+17, 1.297991048295708e+17, 1.297991048336333e+17, 1.297991048376957e+17, 1.29799104841602e+17, 1.297991048456645e+17, 1.29799104849727e+17, 1.297991048536332e+17, 1.297991048576957e+17, 1.297991048617582e+17, 1.297991048658207e+17, 1.29799104869727e+17, 1.297991048737896e+17, 1.29799104877852e+17, 1.297991048817583e+17, 1.297991048858207e+17, 1.297991048898833e+17, 1.297991048937894e+17, 1.297991048978519e+17, 1.297991049019145e+17, 1.297991049058207e+17, 1.297991049098833e+17, 1.297991049139459e+17, 1.297991049180082e+17, 1.297991049219145e+17, 1.29799104925977e+17, 1.297991049300394e+17, 1.297991049339457e+17, 1.297991049380082e+17, 1.297991049420708e+17, 1.297991049461332e+17, 1.297991049500396e+17, 1.29799104954102e+17, 1.297991049581645e+17, 1.297991049620708e+17, 1.297991049661332e+17, 1.297991049701957e+17, 1.29799104974102e+17, 1.297991049781645e+17, 1.297991049822269e+17, 1.297991049862895e+17, 1.297991049901957e+17, 1.297991049942583e+17, 1.297991049983208e+17, 1.297991050022269e+17, 1.297991050062895e+17, 1.29799105010352e+17, 1.297991050144145e+17, 1.297991050183208e+17, 1.297991050223832e+17, 1.297991050264457e+17, 1.29799105030352e+17, 1.297991050344145e+17, 1.297991050384771e+17, 1.297991050423832e+17, 1.297991050464458e+17, 1.297991050505083e+17, 1.297991050545708e+17, 1.297991050584771e+17, 1.297991050625394e+17, 1.29799105066602e+17, 1.297991050705082e+17, 1.297991050745708e+17, 1.297991050786333e+17, 1.297991050825395e+17, 1.29799105086602e+17, 1.297991050906646e+17, 1.297991050945708e+17, 1.297991050986332e+17, 1.297991051026957e+17, 1.297991051067583e+17, 1.297991051106644e+17, 1.29799105114727e+17, 1.297991051187895e+17, 1.297991051226957e+17, 1.297991051267583e+17, 1.297991051308207e+17, 1.297991051348832e+17, 1.297991051387895e+17, 1.29799105142852e+17, 1.297991051469144e+17, 1.297991051508207e+17, 1.297991051548832e+17, 1.297991051589458e+17, 1.29799105162852e+17, 1.297991051669144e+17, 1.29799105170977e+17, 1.297991051750395e+17, 1.297991051789458e+17, 1.297991051830083e+17, 1.297991051870707e+17, 1.29799105190977e+17, 1.297991051950395e+17, 1.29799105199102e+17, 1.297991052031645e+17, 1.297991052070707e+17, 1.297991052111333e+17, 1.297991052151958e+17, 1.297991052191021e+17, 1.297991052231645e+17, 1.297991052272269e+17, 1.297991052311333e+17, 1.297991052351958e+17, 1.297991052392582e+17, 1.297991052433208e+17, 1.29799105247227e+17, 1.297991052512895e+17, 1.297991052553521e+17, 1.297991052592582e+17, 1.297991052633207e+17, 1.297991052673833e+17, 1.297991052712895e+17, 1.297991052753521e+17, 1.297991052794145e+17, 1.297991052833208e+17, 1.297991052873832e+17, 1.297991052914458e+17, 1.297991052955082e+17, 1.297991052994144e+17, 1.29799105303477e+17, 1.297991053075396e+17, 1.297991053114458e+17, 1.297991053155084e+17, 1.297991053195707e+17, 1.297991053236333e+17, 1.297991053275395e+17, 1.297991053316019e+17, 1.297991053356645e+17, 1.297991053395707e+17, 1.297991053436333e+17, 1.297991053476959e+17, 1.29799105351602e+17, 1.297991053556645e+17, 1.29799105359727e+17, 1.297991053637894e+17, 1.297991053676957e+17, 1.297991053717582e+17, 1.297991053758208e+17, 1.29799105379727e+17, 1.297991053837896e+17, 1.29799105387852e+17, 1.297991053919145e+17, 1.297991053958208e+17, 1.297991053998833e+17, 1.297991054039457e+17, 1.29799105407852e+17, 1.297991054119145e+17, 1.29799105415977e+17, 1.297991054198833e+17, 1.297991054239457e+17, 1.297991054280082e+17, 1.297991054320708e+17, 1.29799105435977e+17, 1.297991054400396e+17, 1.29799105444102e+17, 1.297991054480083e+17, 1.297991054520708e+17, 1.297991054561332e+17, 1.297991054600396e+17, 1.297991054641019e+17, 1.297991054681645e+17, 1.297991054720707e+17, 1.297991054761332e+17, 1.297991054801958e+17, 1.297991054842582e+17, 1.297991054881645e+17, 1.297991054922271e+17, 1.297991054962894e+17, 1.297991055001957e+17, 1.297991055042582e+17, 1.297991055083208e+17, 1.297991055123834e+17, 1.297991055162895e+17, 1.29799105520352e+17, 1.297991055244146e+17, 1.297991055283208e+17, 1.297991055323832e+17, 1.297991055364457e+17, 1.29799105540352e+17, 1.297991055444145e+17, 1.297991055484771e+17, 1.297991055525395e+17, 1.297991055564457e+17, 1.297991055605083e+17, 1.297991055645708e+17, 1.297991055684769e+17, 1.297991055725395e+17, 1.29799105576602e+17, 1.297991055806644e+17, 1.297991055845708e+17, 1.297991055886332e+17, 1.297991055926957e+17, 1.29799105596602e+17, 1.297991056006644e+17, 1.29799105604727e+17, 1.297991056086332e+17, 1.297991056126958e+17, 1.297991056167583e+17, 1.297991056208207e+17, 1.29799105624727e+17, 1.297991056287894e+17, 1.29799105632852e+17, 1.297991056367583e+17, 1.297991056408207e+17, 1.297991056448833e+17, 1.297991056487895e+17, 1.29799105652852e+17, 1.297991056569146e+17, 1.297991056608207e+17, 1.297991056648832e+17, 1.297991056689458e+17, 1.297991056730083e+17, 1.297991056769146e+17, 1.29799105680977e+17, 1.297991056850395e+17, 1.297991056889457e+17, 1.297991056930083e+17, 1.297991056970707e+17, 1.297991057011332e+17, 1.297991057050395e+17, 1.297991057091021e+17, 1.297991057131645e+17, 1.297991057170708e+17, 1.297991057211332e+17, 1.297991057251958e+17, 1.29799105729102e+17, 1.297991057331644e+17, 1.29799105737227e+17, 1.297991057412895e+17, 1.297991057451958e+17, 1.297991057492584e+17, 1.297991057533207e+17, 1.29799105757227e+17, 1.297991057612895e+17, 1.297991057653519e+17, 1.297991057694145e+17, 1.297991057733207e+17, 1.297991057773833e+17, 1.297991057814458e+17, 1.297991057853521e+17, 1.297991057894145e+17, 1.29799105793477e+17, 1.297991057973833e+17, 1.297991058014458e+17, 1.297991058055082e+17, 1.297991058095708e+17, 1.29799105813477e+17, 1.297991058175395e+17, 1.29799105821602e+17, 1.297991058255082e+17, 1.297991058295708e+17, 1.297991058336333e+17, 1.297991058375395e+17, 1.29799105841602e+17, 1.297991058456645e+17, 1.297991058495708e+17, 1.297991058536333e+17, 1.297991058576957e+17, 1.297991058617582e+17, 1.297991058656645e+17, 1.29799105869727e+17, 1.297991058737896e+17, 1.297991058776957e+17, 1.297991058817583e+17, 1.297991058858207e+17, 1.297991058898833e+17, 1.297991058937896e+17, 1.297991058978519e+17, 1.297991059019145e+17, 1.297991059058207e+17, 1.297991059098833e+17, 1.297991059139459e+17, 1.29799105917852e+17, 1.297991059219145e+17, 1.297991059259771e+17, 1.297991059300394e+17, 1.297991059339457e+17, 1.297991059380082e+17, 1.297991059420708e+17, 1.29799105945977e+17, 1.297991059500396e+17, 1.29799105954102e+17, 1.297991059581645e+17, 1.297991059620708e+17, 1.297991059661332e+17, 1.297991059701957e+17, 1.29799105974102e+17, 1.297991059781645e+17, 1.297991059822269e+17, 1.297991059861332e+17, 1.297991059901957e+17, 1.297991059942583e+17, 1.297991059983208e+17, 1.297991060022269e+17, 1.297991060062895e+17, 1.29799106010352e+17, 1.297991060142583e+17, 1.297991060183208e+17, 1.297991060223832e+17, 1.297991060262895e+17, 1.29799106030352e+17, 1.297991060344145e+17, 1.297991060383208e+17, 1.297991060423832e+17, 1.297991060464458e+17, 1.297991060505083e+17, 1.297991060544145e+17, 1.297991060584771e+17, 1.297991060625394e+17, 1.297991060664458e+17, 1.297991060705083e+17, 1.297991060745708e+17, 1.297991060786333e+17, 1.297991060825395e+17, 1.29799106086602e+17, 1.297991060906646e+17, 1.297991060945708e+17, 1.297991060986332e+17, 1.297991061026957e+17, 1.29799106106602e+17, 1.297991061106646e+17, 1.29799106114727e+17, 1.297991061187895e+17, 1.297991061226957e+17, 1.297991061267583e+17, 1.297991061308207e+17, 1.297991061347269e+17, 1.297991061387895e+17, 1.29799106142852e+17, 1.297991061469144e+17, 1.297991061508209e+17, 1.297991061548832e+17, 1.297991061589458e+17, 1.29799106162852e+17, 1.297991061669144e+17, 1.29799106170977e+17, 1.297991061748832e+17, 1.297991061789458e+17, 1.297991061830083e+17, 1.297991061870707e+17, 1.29799106190977e+17, 1.297991061950395e+17, 1.29799106199102e+17, 1.297991062030083e+17, 1.297991062070707e+17, 1.297991062111333e+17, 1.297991062150395e+17, 1.29799106219102e+17, 1.297991062231645e+17, 1.297991062270707e+17, 1.297991062311333e+17, 1.297991062351958e+17, 1.297991062392582e+17, 1.297991062431645e+17, 1.29799106247227e+17, 1.297991062512895e+17, 1.297991062551958e+17, 1.297991062592582e+17, 1.297991062633207e+17, 1.297991062673833e+17, 1.297991062712895e+17, 1.297991062753521e+17, 1.297991062794145e+17, 1.297991062833208e+17, 1.297991062873833e+17, 1.297991062914458e+17, 1.297991062953521e+17, 1.297991062994144e+17, 1.29799106303477e+17, 1.297991063075396e+17, 1.297991063114458e+17, 1.297991063155084e+17, 1.297991063195707e+17, 1.29799106323477e+17, 1.297991063275396e+17, 1.297991063316019e+17, 1.297991063356645e+17, 1.297991063395707e+17, 1.297991063436333e+17, 1.297991063476957e+17, 1.29799106351602e+17, 1.297991063556645e+17, 1.29799106359727e+17, 1.297991063636333e+17, 1.297991063676957e+17, 1.297991063717582e+17, 1.297991063758208e+17, 1.29799106379727e+17, 1.297991063837894e+17, 1.29799106387852e+17, 1.297991063917582e+17, 1.297991063958208e+17, 1.297991063998833e+17, 1.297991064037894e+17, 1.29799106407852e+17, 1.297991064119145e+17, 1.297991064158208e+17, 1.297991064198833e+17, 1.297991064239457e+17, 1.297991064280082e+17, 1.297991064319145e+17, 1.29799106435977e+17, 1.297991064400396e+17, 1.297991064439457e+17, 1.297991064480083e+17, 1.297991064520708e+17, 1.297991064561332e+17, 1.297991064600396e+17, 1.297991064641019e+17, 1.297991064681645e+17, 1.297991064720708e+17, 1.297991064761332e+17, 1.297991064801958e+17, 1.29799106484102e+17, 1.297991064881645e+17, 1.297991064922271e+17, 1.297991064962894e+17, 1.297991065001957e+17, 1.297991065042582e+17, 1.297991065083208e+17, 1.297991065122271e+17, 1.297991065162895e+17, 1.29799106520352e+17, 1.297991065244146e+17, 1.297991065283208e+17, 1.297991065323832e+17, 1.297991065364457e+17, 1.29799106540352e+17, 1.297991065444145e+17, 1.297991065484769e+17, 1.297991065523834e+17, 1.297991065564457e+17, 1.297991065605083e+17, 1.297991065645708e+17, 1.297991065684769e+17, 1.297991065725395e+17, 1.29799106576602e+17, 1.297991065805083e+17, 1.297991065845708e+17, 1.297991065886332e+17, 1.297991065925395e+17, 1.29799106596602e+17, 1.297991066006644e+17, 1.297991066045708e+17, 1.297991066086332e+17, 1.297991066126958e+17, 1.297991066167583e+17, 1.297991066206644e+17, 1.29799106624727e+17, 1.297991066287895e+17, 1.297991066326958e+17, 1.297991066367583e+17, 1.297991066408207e+17, 1.297991066448833e+17, 1.297991066487895e+17, 1.29799106652852e+17, 1.297991066569146e+17, 1.297991066608207e+17, 1.297991066648832e+17, 1.297991066689458e+17, 1.29799106672852e+17, 1.297991066769146e+17, 1.29799106680977e+17, 1.297991066850395e+17, 1.297991066889458e+17, 1.297991066930083e+17, 1.297991066970707e+17, 1.297991067009769e+17, 1.297991067050395e+17, 1.297991067091021e+17, 1.297991067131644e+17, 1.297991067170708e+17, 1.297991067211332e+17, 1.297991067251958e+17, 1.297991067291021e+17, 1.297991067331644e+17, 1.29799106737227e+17, 1.297991067411332e+17, 1.297991067451958e+17, 1.297991067492582e+17, 1.297991067533207e+17, 1.29799106757227e+17, 1.297991067612895e+17, 1.297991067653519e+17, 1.297991067692582e+17, 1.297991067733207e+17, 1.297991067773833e+17, 1.297991067812895e+17, 1.297991067853519e+17, 1.297991067894145e+17, 1.297991067933207e+17, 1.297991067973833e+17, 1.297991068014458e+17, 1.297991068055082e+17, 1.297991068094145e+17, 1.29799106813477e+17, 1.297991068175395e+17, 1.297991068214458e+17, 1.297991068255082e+17, 1.297991068295707e+17, 1.297991068336333e+17, 1.297991068375395e+17, 1.29799106841602e+17, 1.297991068456645e+17, 1.297991068495708e+17, 1.297991068536333e+17, 1.297991068576957e+17, 1.29799106861602e+17, 1.297991068656644e+17, 1.29799106869727e+17, 1.297991068737896e+17, 1.297991068776957e+17, 1.297991068817583e+17, 1.297991068858208e+17, 1.29799106889727e+17, 1.297991068937896e+17, 1.297991068978519e+17, 1.297991069019145e+17, 1.297991069058207e+17, 1.297991069098833e+17, 1.297991069139457e+17, 1.29799106917852e+17, 1.297991069219145e+17, 1.297991069259771e+17, 1.297991069298833e+17, 1.297991069339457e+17, 1.297991069380082e+17, 1.297991069420708e+17, 1.297991069459771e+17, 1.297991069500394e+17, 1.29799106954102e+17, 1.297991069580082e+17, 1.297991069620708e+17, 1.297991069661332e+17, 1.297991069700394e+17, 1.29799106974102e+17, 1.297991069781645e+17, 1.297991069820708e+17, 1.297991069861332e+17, 1.297991069901957e+17, 1.297991069942582e+17, 1.297991069981645e+17, 1.297991070022269e+17, 1.297991070062895e+17, 1.297991070101957e+17, 1.297991070142583e+17, 1.297991070183208e+17, 1.297991070223832e+17, 1.297991070262895e+17, 1.29799107030352e+17, 1.297991070344145e+17, 1.297991070383208e+17, 1.297991070423832e+17, 1.297991070464458e+17, 1.29799107050352e+17, 1.297991070544145e+17, 1.297991070584771e+17, 1.297991070625395e+17, 1.297991070664457e+17, 1.297991070705083e+17, 1.297991070745708e+17, 1.297991070784771e+17, 1.297991070825395e+17, 1.29799107086602e+17, 1.297991070906646e+17, 1.297991070945708e+17, 1.297991070986332e+17, 1.297991071026958e+17, 1.29799107106602e+17, 1.297991071106646e+17, 1.297991071147269e+17, 1.297991071186333e+17, 1.297991071226957e+17, 1.297991071267583e+17, 1.297991071308207e+17, 1.297991071347269e+17, 1.297991071387895e+17, 1.297991071428521e+17, 1.297991071467583e+17, 1.297991071508207e+17, 1.297991071548832e+17, 1.297991071587895e+17, 1.29799107162852e+17, 1.297991071669144e+17, 1.297991071708207e+17, 1.297991071748832e+17, 1.297991071789458e+17, 1.297991071830083e+17, 1.297991071869146e+17, 1.29799107190977e+17, 1.297991071950395e+17, 1.297991071989458e+17, 1.297991072030083e+17, 1.297991072070707e+17, 1.297991072111333e+17, 1.297991072150395e+17, 1.29799107219102e+17, 1.297991072231645e+17, 1.297991072270707e+17, 1.297991072311332e+17, 1.297991072351958e+17, 1.29799107239102e+17, 1.297991072431645e+17, 1.29799107247227e+17, 1.297991072512895e+17, 1.297991072551958e+17, 1.297991072592582e+17, 1.297991072633207e+17, 1.297991072672269e+17, 1.297991072712895e+17, 1.297991072753521e+17, 1.297991072794144e+17, 1.297991072833208e+17, 1.297991072873833e+17, 1.297991072914458e+17, 1.297991072953521e+17, 1.297991072994144e+17, 1.29799107303477e+17, 1.297991073073832e+17, 1.297991073114458e+17, 1.297991073155084e+17, 1.297991073195708e+17, 1.29799107323477e+17, 1.297991073275396e+17, 1.297991073316019e+17, 1.297991073355082e+17, 1.297991073395707e+17, 1.297991073436333e+17, 1.297991073475396e+17, 1.29799107351602e+17, 1.297991073556645e+17, 1.297991073595707e+17, 1.297991073636333e+17, 1.297991073676957e+17, 1.297991073717582e+17, 1.297991073756645e+17, 1.29799107379727e+17, 1.297991073837894e+17, 1.297991073876959e+17, 1.297991073917582e+17, 1.297991073958207e+17, 1.297991073998833e+17, 1.297991074037894e+17, 1.29799107407852e+17, 1.297991074119145e+17, 1.297991074158208e+17, 1.297991074198833e+17, 1.297991074239457e+17, 1.29799107427852e+17, 1.297991074319145e+17, 1.29799107435977e+17, 1.297991074400396e+17, 1.297991074439457e+17, 1.297991074480083e+17, 1.297991074520708e+17, 1.29799107455977e+17, 1.297991074600396e+17, 1.29799107464102e+17, 1.297991074681645e+17, 1.297991074720708e+17, 1.297991074761332e+17, 1.297991074801958e+17, 1.29799107484102e+17, 1.297991074881645e+17, 1.297991074922271e+17, 1.297991074961332e+17, 1.297991075001957e+17, 1.297991075042583e+17, 1.297991075083208e+17, 1.297991075122271e+17, 1.297991075162895e+17, 1.29799107520352e+17, 1.297991075242582e+17, 1.297991075283208e+17, 1.297991075323832e+17, 1.297991075362894e+17, 1.29799107540352e+17, 1.297991075444146e+17, 1.297991075483208e+17, 1.297991075523834e+17, 1.297991075564457e+17, 1.297991075605082e+17, 1.297991075644145e+17, 1.297991075684769e+17, 1.297991075725395e+17, 1.297991075764457e+17, 1.297991075805083e+17, 1.297991075845708e+17, 1.297991075886332e+17, 1.297991075925395e+17, 1.29799107596602e+17, 1.297991076006644e+17, 1.297991076045708e+17, 1.297991076086332e+17, 1.297991076126958e+17, 1.29799107616602e+17, 1.297991076206644e+17, 1.29799107624727e+17, 1.297991076287895e+17, 1.297991076326957e+17, 1.297991076367583e+17, 1.297991076408207e+17, 1.29799107644727e+17, 1.297991076487895e+17, 1.29799107652852e+17, 1.297991076569146e+17, 1.297991076608207e+17, 1.297991076648832e+17, 1.297991076689458e+17, 1.29799107672852e+17, 1.297991076769146e+17, 1.29799107680977e+17, 1.297991076848833e+17, 1.297991076889458e+17, 1.297991076930083e+17, 1.297991076970707e+17, 1.297991077009769e+17, 1.297991077050395e+17, 1.297991077091021e+17, 1.297991077130083e+17, 1.297991077170708e+17, 1.297991077211333e+17, 1.297991077250395e+17, 1.297991077291021e+17, 1.297991077331644e+17, 1.297991077370707e+17, 1.297991077411332e+17, 1.297991077451958e+17, 1.297991077492582e+17, 1.297991077531645e+17, 1.29799107757227e+17, 1.297991077612895e+17, 1.297991077651958e+17, 1.297991077692582e+17, 1.297991077733207e+17, 1.297991077773833e+17, 1.297991077812895e+17, 1.297991077853519e+17, 1.297991077894145e+17, 1.297991077933207e+17, 1.297991077973832e+17, 1.297991078014458e+17, 1.297991078053519e+17, 1.297991078094145e+17, 1.29799107813477e+17, 1.297991078175395e+17, 1.297991078214458e+17, 1.297991078255082e+17, 1.297991078295707e+17, 1.29799107833477e+17, 1.297991078375395e+17, 1.29799107841602e+17, 1.297991078456645e+17, 1.297991078495708e+17, 1.297991078536333e+17, 1.297991078576957e+17, 1.29799107861602e+17, 1.297991078656645e+17, 1.29799107869727e+17, 1.297991078736333e+17, 1.297991078776957e+17, 1.297991078817583e+17, 1.297991078858208e+17, 1.29799107889727e+17, 1.297991078937896e+17, 1.297991078978519e+17, 1.297991079017582e+17, 1.297991079058208e+17, 1.297991079098833e+17, 1.297991079137896e+17, 1.29799107917852e+17, 1.297991079219145e+17, 1.297991079258207e+17, 1.297991079298833e+17, 1.297991079339457e+17, 1.297991079380083e+17, 1.297991079419145e+17, 1.297991079459771e+17, 1.297991079500394e+17, 1.297991079539459e+17, 1.297991079580082e+17, 1.297991079620707e+17, 1.297991079661332e+17, 1.297991079700394e+17, 1.29799107974102e+17, 1.297991079781646e+17, 1.297991079820708e+17, 1.297991079861332e+17, 1.297991079901957e+17, 1.29799107994102e+17, 1.297991079981645e+17, 1.297991080022269e+17, 1.297991080062895e+17, 1.297991080101957e+17, 1.297991080142583e+17, 1.297991080183208e+17, 1.297991080222269e+17, 1.297991080262895e+17, 1.29799108030352e+17, 1.297991080344145e+17, 1.297991080383208e+17, 1.297991080423832e+17, 1.297991080464458e+17, 1.29799108050352e+17, 1.297991080544145e+17, 1.297991080584771e+17, 1.297991080623832e+17, 1.297991080664457e+17, 1.297991080705083e+17, 1.297991080745708e+17, 1.297991080784771e+17, 1.297991080825395e+17, 1.29799108086602e+17, 1.297991080905083e+17, 1.297991080945708e+17, 1.297991080986332e+17, 1.297991081025394e+17, 1.29799108106602e+17, 1.297991081106646e+17, 1.297991081145708e+17, 1.297991081186333e+17, 1.297991081226958e+17, 1.297991081267583e+17, 1.297991081306646e+17, 1.297991081347269e+17, 1.297991081387895e+17, 1.297991081426957e+17, 1.297991081467583e+17, 1.297991081508207e+17, 1.297991081548832e+17, 1.297991081587895e+17, 1.297991081628521e+17, 1.297991081669144e+17, 1.297991081708207e+17, 1.297991081748832e+17, 1.297991081789458e+17, 1.29799108182852e+17, 1.297991081869144e+17, 1.29799108190977e+17, 1.297991081950395e+17, 1.297991081989458e+17, 1.297991082030083e+17, 1.297991082070707e+17, 1.29799108210977e+17, 1.297991082150395e+17, 1.29799108219102e+17, 1.297991082231645e+17, 1.297991082270707e+17, 1.297991082311332e+17, 1.297991082351958e+17, 1.29799108239102e+17, 1.297991082431645e+17, 1.29799108247227e+17, 1.297991082511333e+17, 1.297991082551958e+17, 1.297991082592582e+17, 1.297991082633207e+17, 1.29799108267227e+17, 1.297991082712895e+17, 1.297991082753521e+17, 1.297991082792582e+17, 1.297991082833208e+17, 1.297991082873833e+17, 1.297991082912895e+17, 1.297991082953521e+17, 1.297991082994144e+17, 1.297991083033207e+17, 1.297991083073833e+17, 1.297991083114458e+17, 1.297991083155082e+17, 1.297991083194145e+17, 1.29799108323477e+17, 1.297991083275396e+17, 1.297991083314458e+17, 1.297991083355082e+17, 1.297991083395708e+17, 1.297991083436333e+17, 1.297991083475396e+17, 1.297991083516019e+17, 1.297991083556645e+17, 1.297991083595707e+17, 1.297991083636333e+17, 1.297991083676957e+17, 1.297991083716019e+17, 1.297991083756645e+17, 1.297991083797271e+17, 1.297991083837894e+17, 1.297991083876957e+17, 1.297991083917582e+17, 1.297991083958207e+17, 1.29799108399727e+17, 1.297991084037894e+17, 1.29799108407852e+17, 1.297991084119145e+17, 1.297991084158208e+17, 1.297991084198833e+17, 1.297991084239457e+17, 1.29799108427852e+17, 1.297991084319145e+17, 1.29799108435977e+17, 1.297991084398833e+17, 1.297991084439457e+17, 1.297991084480083e+17, 1.297991084520708e+17, 1.29799108455977e+17, 1.297991084600396e+17, 1.29799108464102e+17, 1.297991084680082e+17, 1.297991084720708e+17, 1.297991084761332e+17, 1.297991084800396e+17, 1.29799108484102e+17, 1.297991084881645e+17, 1.297991084920708e+17, 1.297991084961332e+17, 1.297991085001957e+17, 1.297991085042583e+17, 1.297991085081645e+17, 1.297991085122271e+17, 1.297991085162894e+17, 1.297991085201958e+17, 1.297991085242583e+17, 1.297991085283208e+17, 1.297991085323832e+17, 1.297991085362894e+17, 1.29799108540352e+17, 1.297991085444146e+17, 1.297991085483208e+17, 1.297991085523832e+17, 1.297991085564457e+17, 1.29799108560352e+17, 1.297991085644146e+17, 1.297991085684769e+17, 1.297991085725395e+17, 1.297991085764457e+17, 1.297991085805083e+17, 1.297991085845708e+17, 1.297991085884769e+17, 1.297991085925395e+17, 1.29799108596602e+17, 1.297991086006644e+17, 1.297991086045708e+17, 1.297991086086332e+17, 1.297991086126958e+17, 1.29799108616602e+17, 1.297991086206644e+17, 1.29799108624727e+17, 1.297991086286332e+17, 1.297991086326957e+17, 1.297991086367583e+17, 1.297991086408207e+17, 1.29799108644727e+17, 1.297991086487895e+17, 1.29799108652852e+17, 1.297991086567583e+17, 1.297991086608207e+17, 1.297991086648832e+17, 1.297991086687895e+17, 1.29799108672852e+17, 1.297991086769146e+17, 1.297991086808207e+17, 1.297991086848833e+17, 1.297991086889458e+17, 1.297991086930083e+17, 1.297991086969146e+17, 1.29799108700977e+17, 1.297991087050395e+17, 1.297991087089458e+17, 1.297991087130083e+17, 1.297991087170707e+17, 1.297991087211333e+17, 1.297991087250395e+17, 1.297991087291021e+17, 1.297991087331644e+17, 1.297991087370707e+17, 1.297991087411333e+17, 1.297991087451958e+17, 1.297991087491021e+17, 1.297991087531644e+17, 1.29799108757227e+17, 1.297991087612895e+17, 1.297991087651958e+17, 1.297991087692582e+17, 1.297991087733207e+17, 1.29799108777227e+17, 1.297991087812896e+17, 1.297991087853519e+17, 1.297991087894145e+17, 1.297991087933207e+17, 1.297991087973832e+17, 1.297991088014458e+17, 1.297991088053519e+17, 1.297991088094145e+17, 1.29799108813477e+17, 1.297991088173833e+17, 1.297991088214458e+17, 1.297991088255082e+17, 1.297991088295707e+17, 1.29799108833477e+17, 1.297991088375395e+17, 1.29799108841602e+17, 1.297991088455082e+17, 1.297991088495708e+17, 1.297991088536333e+17, 1.297991088575395e+17, 1.29799108861602e+17, 1.297991088656645e+17, 1.297991088695707e+17, 1.297991088736333e+17, 1.297991088776957e+17, 1.297991088817582e+17, 1.297991088856645e+17, 1.29799108889727e+17, 1.297991088937896e+17, 1.297991088976957e+17, 1.297991089017582e+17, 1.297991089058208e+17, 1.297991089098833e+17, 1.297991089137896e+17, 1.297991089178519e+17, 1.297991089219145e+17, 1.297991089258208e+17, 1.297991089298833e+17, 1.297991089339457e+17, 1.297991089378519e+17, 1.297991089419145e+17, 1.297991089459771e+17, 1.297991089500394e+17, 1.297991089539457e+17, 1.297991089580082e+17, 1.297991089620707e+17, 1.297991089659771e+17, 1.297991089700394e+17, 1.29799108974102e+17, 1.297991089781646e+17, 1.297991089820708e+17, 1.297991089861332e+17, 1.297991089901957e+17, 1.29799108994102e+17, 1.297991089981645e+17, 1.297991090022269e+17, 1.297991090061332e+17, 1.297991090101957e+17, 1.297991090142583e+17, 1.297991090183208e+17, 1.297991090222269e+17, 1.297991090262895e+17, 1.29799109030352e+17, 1.297991090342582e+17, 1.297991090383208e+17, 1.297991090423832e+17, 1.297991090462895e+17, 1.29799109050352e+17, 1.297991090544145e+17, 1.297991090583208e+17, 1.297991090623832e+17, 1.297991090664457e+17, 1.297991090705083e+17, 1.297991090744145e+17, 1.297991090784771e+17, 1.297991090825395e+17, 1.297991090864458e+17, 1.297991090905083e+17, 1.297991090945708e+17, 1.297991090986332e+17, 1.297991091025395e+17, 1.29799109106602e+17, 1.297991091106646e+17, 1.297991091145708e+17, 1.297991091186332e+17, 1.297991091226958e+17, 1.29799109126602e+17, 1.297991091306646e+17, 1.297991091347269e+17, 1.297991091387895e+17, 1.297991091426958e+17, 1.297991091467583e+17, 1.297991091508207e+17, 1.297991091547269e+17, 1.297991091587895e+17, 1.29799109162852e+17, 1.297991091669144e+17, 1.297991091708207e+17, 1.297991091748832e+17, 1.297991091789458e+17, 1.297991091828521e+17, 1.297991091869144e+17, 1.29799109190977e+17, 1.297991091948832e+17, 1.297991091989457e+17, 1.297991092030083e+17, 1.297991092070707e+17, 1.29799109210977e+17, 1.297991092150395e+17, 1.29799109219102e+17, 1.297991092230083e+17, 1.297991092270707e+17, 1.297991092311332e+17, 1.297991092350395e+17, 1.29799109239102e+17, 1.297991092431645e+17, 1.297991092470707e+17, 1.297991092511333e+17, 1.297991092551958e+17, 1.297991092592582e+17, 1.297991092631645e+17, 1.29799109267227e+17, 1.297991092712895e+17, 1.297991092751958e+17, 1.297991092792582e+17, 1.297991092833207e+17, 1.297991092873833e+17, 1.297991092912895e+17, 1.297991092953521e+17, 1.297991092994145e+17, 1.297991093033207e+17, 1.297991093073833e+17, 1.297991093114458e+17, 1.297991093153521e+17, 1.297991093194145e+17, 1.29799109323477e+17, 1.297991093275395e+17, 1.297991093314458e+17, 1.297991093355082e+17, 1.297991093395708e+17, 1.29799109343477e+17, 1.297991093475396e+17, 1.297991093516019e+17, 1.297991093556645e+17, 1.297991093595708e+17, 1.297991093636332e+17, 1.297991093676957e+17, 1.297991093716019e+17, 1.297991093756645e+17, 1.297991093797271e+17, 1.297991093836333e+17, 1.297991093876957e+17, 1.297991093917582e+17, 1.297991093958207e+17, 1.29799109399727e+17, 1.297991094037894e+17, 1.29799109407852e+17, 1.297991094117582e+17, 1.297991094158208e+17, 1.297991094198833e+17, 1.297991094237894e+17, 1.29799109427852e+17, 1.297991094319145e+17, 1.297991094358207e+17, 1.297991094398833e+17, 1.297991094439457e+17, 1.297991094480083e+17, 1.297991094519145e+17, 1.29799109455977e+17, 1.297991094600396e+17, 1.297991094639457e+17, 1.297991094680082e+17, 1.297991094720708e+17, 1.297991094761332e+17, 1.297991094800396e+17, 1.29799109484102e+17, 1.297991094881645e+17, 1.297991094920708e+17, 1.297991094961332e+17, 1.297991095001957e+17, 1.29799109504102e+17, 1.297991095081645e+17, 1.297991095122271e+17, 1.297991095162895e+17, 1.297991095201958e+17, 1.297991095242583e+17, 1.297991095283206e+17, 1.297991095322271e+17, 1.297991095362894e+17, 1.29799109540352e+17, 1.297991095444146e+17, 1.297991095483208e+17, 1.297991095523832e+17, 1.297991095564458e+17, 1.29799109560352e+17, 1.297991095644145e+17, 1.297991095684769e+17, 1.297991095723832e+17, 1.297991095764457e+17, 1.297991095805083e+17, 1.297991095845708e+17, 1.297991095884769e+17, 1.297991095925395e+17, 1.29799109596602e+17, 1.297991096005082e+17, 1.297991096045708e+17, 1.297991096086332e+17, 1.297991096125395e+17, 1.297991096166021e+17, 1.297991096206644e+17, 1.297991096245708e+17, 1.297991096286332e+17, 1.297991096326957e+17, 1.297991096367583e+17, 1.297991096406644e+17, 1.29799109644727e+17, 1.297991096487895e+17, 1.297991096526958e+17, 1.297991096567583e+17, 1.297991096608207e+17, 1.297991096648832e+17, 1.297991096687895e+17, 1.29799109672852e+17, 1.297991096769146e+17, 1.297991096808207e+17, 1.297991096848833e+17, 1.297991096889458e+17, 1.29799109692852e+17, 1.297991096969146e+17, 1.29799109700977e+17, 1.297991097050395e+17, 1.297991097089458e+17, 1.297991097130083e+17, 1.297991097170707e+17, 1.29799109720977e+17, 1.297991097250395e+17, 1.29799109729102e+17, 1.297991097331645e+17, 1.297991097370707e+17, 1.297991097411333e+17, 1.297991097451958e+17, 1.297991097491021e+17, 1.297991097531644e+17, 1.29799109757227e+17, 1.297991097611333e+17, 1.297991097651956e+17, 1.297991097692582e+17, 1.297991097733208e+17, 1.29799109777227e+17, 1.297991097812896e+17, 1.297991097853519e+17, 1.297991097892582e+17, 1.297991097933207e+17, 1.297991097973832e+17, 1.297991098012895e+17, 1.297991098053519e+17, 1.297991098094145e+17, 1.297991098133207e+17, 1.297991098173833e+17, 1.297991098214458e+17, 1.297991098255082e+17, 1.297991098294145e+17, 1.29799109833477e+17, 1.297991098375395e+17, 1.297991098414458e+17, 1.297991098455082e+17, 1.297991098495708e+17, 1.297991098536333e+17, 1.297991098575395e+17, 1.29799109861602e+17, 1.297991098656645e+17, 1.297991098695707e+17, 1.297991098736333e+17, 1.297991098776957e+17, 1.29799109881602e+17, 1.297991098856645e+17, 1.29799109889727e+17, 1.297991098937894e+17, 1.297991098976957e+17, 1.297991099017582e+17, 1.297991099058208e+17, 1.29799109909727e+17, 1.297991099137896e+17, 1.29799109917852e+17, 1.297991099219145e+17, 1.297991099258208e+17, 1.297991099298831e+17, 1.297991099339457e+17, 1.297991099378519e+17, 1.297991099419145e+17, 1.297991099459771e+17, 1.297991099498833e+17, 1.297991099539457e+17, 1.297991099580083e+17, 1.297991099620707e+17, 1.29799109965977e+17, 1.297991099700394e+17, 1.29799109974102e+17, 1.297991099780082e+17, 1.297991099820708e+17, 1.297991099861332e+17, 1.297991099900394e+17, 1.29799109994102e+17, 1.297991099981645e+17, 1.297991100020708e+17, 1.297991100061332e+17, 1.297991100101957e+17, 1.297991100142583e+17, 1.297991100181646e+17, 1.297991100222269e+17, 1.297991100262895e+17, 1.297991100301957e+17, 1.297991100342582e+17, 1.297991100383208e+17, 1.297991100423832e+17, 1.297991100462895e+17, 1.29799110050352e+17, 1.297991100544145e+17, 1.297991100583208e+17, 1.297991100623832e+17, 1.297991100664457e+17, 1.29799110070352e+17, 1.297991100744145e+17, 1.297991100784771e+17, 1.297991100825395e+17, 1.297991100864458e+17, 1.297991100905083e+17, 1.297991100945708e+17, 1.297991100984771e+17, 1.297991101025395e+17, 1.29799110106602e+17, 1.297991101106646e+17, 1.297991101145708e+17, 1.297991101186332e+17, 1.297991101226958e+17, 1.29799110126602e+17, 1.297991101306646e+17, 1.29799110134727e+17, 1.297991101386332e+17, 1.297991101426958e+17, 1.297991101467583e+17, 1.297991101508207e+17, 1.297991101547269e+17, 1.297991101587895e+17, 1.29799110162852e+17, 1.297991101667583e+17, 1.297991101708207e+17, 1.297991101748833e+17, 1.297991101787895e+17, 1.297991101828521e+17, 1.297991101869144e+17, 1.297991101908207e+17, 1.297991101948832e+17, 1.297991101989457e+17, 1.297991102030083e+17, 1.297991102069144e+17, 1.29799110210977e+17, 1.297991102150396e+17, 1.297991102189458e+17, 1.297991102230083e+17, 1.297991102270707e+17, 1.297991102311332e+17, 1.297991102350395e+17, 1.29799110239102e+17, 1.297991102431645e+17, 1.297991102470707e+17, 1.297991102511333e+17, 1.297991102551958e+17, 1.29799110259102e+17, 1.297991102631645e+17, 1.29799110267227e+17, 1.297991102712895e+17, 1.297991102751958e+17, 1.297991102792582e+17, 1.297991102833207e+17, 1.29799110287227e+17, 1.297991102912895e+17, 1.297991102953521e+17, 1.297991102994145e+17, 1.297991103033207e+17, 1.297991103073833e+17, 1.297991103114458e+17, 1.297991103153521e+17, 1.297991103194145e+17, 1.29799110323477e+17, 1.297991103273833e+17, 1.297991103314458e+17, 1.297991103355082e+17, 1.297991103395708e+17, 1.29799110343477e+17, 1.297991103475396e+17, 1.29799110351602e+17, 1.297991103555082e+17, 1.297991103595708e+17, 1.297991103636332e+17, 1.297991103675396e+17, 1.297991103716019e+17, 1.297991103756645e+17, 1.297991103795708e+17, 1.297991103836333e+17, 1.297991103876957e+17, 1.297991103917583e+17, 1.297991103956645e+17, 1.29799110399727e+17, 1.297991104037894e+17, 1.297991104076957e+17, 1.297991104117582e+17, 1.297991104158208e+17, 1.297991104198833e+17, 1.297991104237894e+17, 1.29799110427852e+17, 1.297991104319145e+17, 1.297991104358207e+17, 1.297991104398833e+17, 1.297991104439457e+17, 1.29799110447852e+17, 1.297991104519145e+17, 1.29799110455977e+17, 1.297991104600396e+17, 1.297991104639457e+17, 1.297991104680082e+17, 1.297991104720708e+17, 1.29799110475977e+17, 1.297991104800396e+17, 1.29799110484102e+17, 1.297991104881645e+17, 1.297991104920708e+17, 1.297991104961332e+17, 1.297991105001957e+17, 1.29799110504102e+17, 1.297991105081645e+17, 1.297991105122271e+17, 1.297991105161332e+17, 1.297991105201957e+17, 1.297991105242583e+17, 1.297991105283206e+17, 1.297991105322271e+17, 1.297991105362895e+17, 1.29799110540352e+17, 1.297991105442583e+17, 1.297991105483208e+17, 1.297991105523832e+17, 1.297991105562894e+17, 1.29799110560352e+17, 1.297991105644145e+17, 1.297991105683208e+17, 1.297991105723832e+17, 1.297991105764458e+17, 1.297991105805083e+17, 1.297991105844146e+17, 1.297991105884769e+17, 1.297991105925395e+17, 1.297991105964457e+17, 1.297991106005082e+17, 1.297991106045708e+17, 1.297991106086332e+17, 1.297991106125395e+17, 1.297991106166021e+17, 1.297991106206644e+17, 1.297991106245708e+17, 1.297991106286332e+17, 1.297991106326957e+17, 1.29799110636602e+17, 1.297991106406644e+17, 1.29799110644727e+17, 1.297991106487895e+17, 1.297991106526958e+17, 1.297991106567583e+17, 1.297991106608207e+17, 1.29799110664727e+17, 1.297991106687895e+17, 1.29799110672852e+17, 1.297991106769146e+17, 1.297991106808207e+17, 1.297991106848832e+17, 1.297991106889458e+17, 1.29799110692852e+17, 1.297991106969146e+17, 1.29799110700977e+17, 1.297991107048832e+17, 1.297991107089458e+17, 1.297991107130083e+17, 1.297991107170707e+17, 1.29799110720977e+17, 1.297991107250395e+17, 1.29799110729102e+17, 1.297991107330083e+17, 1.297991107370707e+17, 1.297991107411333e+17, 1.297991107450395e+17, 1.297991107491021e+17, 1.297991107531645e+17, 1.297991107570707e+17, 1.297991107611333e+17, 1.297991107651956e+17, 1.297991107692582e+17, 1.297991107731644e+17, 1.29799110777227e+17, 1.297991107812896e+17, 1.297991107851958e+17, 1.297991107892582e+17, 1.297991107933208e+17, 1.297991107973832e+17, 1.297991108012895e+17, 1.297991108053519e+17, 1.297991108094145e+17, 1.297991108133207e+17, 1.297991108173833e+17, 1.297991108214458e+17, 1.297991108253519e+17, 1.297991108294145e+17, 1.29799110833477e+17, 1.297991108375395e+17, 1.297991108414458e+17, 1.297991108455082e+17, 1.297991108495707e+17, 1.29799110853477e+17, 1.297991108575395e+17, 1.29799110861602e+17, 1.297991108656645e+17, 1.297991108695707e+17, 1.297991108736333e+17, 1.297991108776957e+17, 1.29799110881602e+17, 1.297991108856645e+17, 1.29799110889727e+17, 1.297991108936333e+17, 1.297991108976957e+17, 1.297991109017582e+17, 1.297991109058208e+17, 1.29799110909727e+17, 1.297991109137896e+17, 1.29799110917852e+17, 1.297991109217582e+17, 1.297991109258208e+17, 1.297991109298831e+17, 1.297991109337896e+17, 1.29799110937852e+17, 1.297991109419145e+17, 1.297991109458208e+17, 1.297991109498833e+17, 1.297991109539457e+17, 1.297991109580083e+17, 1.297991109619145e+17, 1.29799110965977e+17, 1.297991109700394e+17, 1.297991109739457e+17, 1.297991109780083e+17, 1.297991109820708e+17, 1.297991109861332e+17, 1.297991109900394e+17, 1.29799110994102e+17, 1.297991109981645e+17, 1.297991110020707e+17, 1.297991110061332e+17, 1.297991110101958e+17, 1.29799111014102e+17, 1.297991110181646e+17, 1.297991110222269e+17, 1.297991110262895e+17, 1.297991110301957e+17, 1.297991110342582e+17, 1.297991110383208e+17, 1.297991110422269e+17, 1.297991110462895e+17, 1.29799111050352e+17, 1.297991110544145e+17, 1.297991110583208e+17, 1.297991110623832e+17, 1.297991110664457e+17, 1.29799111070352e+17, 1.297991110744145e+17, 1.297991110784771e+17, 1.297991110823832e+17, 1.297991110864457e+17, 1.297991110905083e+17, 1.297991110945708e+17, 1.297991110984771e+17, 1.297991111025395e+17, 1.29799111106602e+17, 1.297991111105083e+17, 1.297991111145708e+17, 1.297991111186332e+17, 1.297991111225395e+17, 1.29799111126602e+17, 1.297991111306644e+17, 1.297991111345708e+17, 1.297991111386332e+17, 1.297991111426958e+17, 1.297991111467583e+17, 1.297991111506646e+17, 1.29799111154727e+17, 1.297991111587895e+17, 1.297991111626958e+17, 1.297991111667581e+17, 1.297991111708207e+17, 1.297991111748833e+17, 1.297991111787895e+17, 1.297991111828521e+17, 1.297991111869144e+17, 1.297991111908207e+17, 1.297991111948833e+17, 1.297991111989457e+17, 1.29799111202852e+17, 1.297991112069144e+17, 1.29799111210977e+17, 1.297991112150395e+17, 1.297991112189458e+17, 1.297991112230083e+17, 1.297991112270707e+17, 1.29799111230977e+17, 1.297991112350395e+17, 1.29799111239102e+17, 1.297991112431645e+17, 1.297991112470707e+17, 1.297991112511332e+17, 1.297991112551958e+17, 1.29799111259102e+17, 1.297991112631645e+17, 1.29799111267227e+17, 1.297991112711332e+17, 1.297991112751958e+17, 1.297991112792582e+17, 1.297991112833207e+17, 1.29799111287227e+17, 1.297991112912895e+17, 1.297991112953519e+17, 1.297991112992582e+17, 1.297991113033207e+17, 1.297991113073833e+17, 1.297991113112895e+17, 1.297991113153521e+17, 1.297991113194145e+17, 1.297991113233208e+17, 1.297991113273833e+17, 1.297991113314456e+17, 1.297991113355082e+17, 1.297991113394145e+17, 1.29799111343477e+17, 1.297991113475396e+17, 1.297991113514458e+17, 1.297991113555082e+17, 1.297991113595708e+17, 1.297991113636332e+17, 1.297991113675395e+17, 1.297991113716019e+17, 1.297991113756645e+17, 1.297991113795708e+17, 1.297991113836333e+17, 1.297991113876957e+17, 1.297991113916019e+17, 1.297991113956645e+17, 1.29799111399727e+17, 1.297991114037894e+17, 1.297991114076957e+17, 1.297991114117583e+17, 1.297991114158207e+17, 1.297991114197271e+17, 1.297991114237894e+17, 1.29799111427852e+17, 1.297991114319145e+17, 1.297991114358207e+17, 1.297991114398833e+17, 1.297991114439457e+17, 1.29799111447852e+17, 1.297991114519146e+17, 1.29799111455977e+17, 1.297991114598833e+17, 1.297991114639457e+17, 1.297991114680082e+17, 1.297991114720708e+17, 1.29799111475977e+17, 1.297991114800396e+17, 1.29799111484102e+17, 1.297991114880083e+17, 1.297991114920708e+17, 1.297991114961332e+17, 1.297991115000396e+17, 1.29799111504102e+17, 1.297991115081645e+17, 1.297991115120708e+17, 1.297991115161332e+17, 1.297991115201957e+17, 1.297991115242583e+17, 1.297991115281645e+17, 1.297991115322269e+17, 1.297991115362895e+17, 1.297991115401957e+17, 1.297991115442583e+17, 1.297991115483208e+17, 1.297991115523832e+17, 1.297991115562895e+17, 1.29799111560352e+17, 1.297991115644145e+17, 1.297991115683206e+17, 1.297991115723832e+17, 1.297991115764458e+17, 1.29799111580352e+17, 1.297991115844146e+17, 1.297991115884769e+17, 1.297991115925395e+17, 1.297991115964458e+17, 1.297991116005082e+17, 1.297991116045708e+17, 1.297991116084769e+17, 1.297991116125395e+17, 1.297991116166021e+17, 1.297991116206644e+17, 1.297991116245708e+17, 1.297991116286332e+17, 1.297991116326957e+17, 1.29799111636602e+17, 1.297991116406644e+17, 1.29799111644727e+17, 1.297991116486332e+17, 1.297991116526958e+17, 1.297991116567583e+17, 1.297991116608207e+17, 1.29799111664727e+17, 1.297991116687895e+17, 1.29799111672852e+17, 1.297991116767583e+17, 1.297991116808207e+17, 1.297991116848832e+17, 1.297991116887895e+17, 1.29799111692852e+17, 1.297991116969144e+17, 1.297991117008207e+17, 1.297991117048832e+17, 1.297991117089458e+17, 1.297991117130083e+17, 1.297991117169146e+17, 1.29799111720977e+17, 1.297991117250395e+17, 1.297991117289458e+17, 1.297991117330081e+17, 1.297991117370707e+17, 1.297991117411333e+17, 1.297991117450395e+17, 1.297991117491021e+17, 1.297991117531645e+17, 1.297991117570707e+17, 1.297991117611333e+17, 1.297991117651956e+17, 1.29799111769102e+17, 1.297991117731645e+17, 1.29799111777227e+17, 1.297991117812896e+17, 1.297991117851958e+17, 1.297991117892582e+17, 1.297991117933208e+17, 1.29799111797227e+17, 1.297991118012895e+17, 1.297991118053519e+17, 1.297991118094145e+17, 1.297991118133208e+17, 1.297991118173833e+17, 1.297991118214458e+17, 1.297991118253519e+17, 1.297991118294145e+17, 1.29799111833477e+17, 1.297991118373832e+17, 1.297991118414458e+17, 1.297991118455082e+17, 1.297991118495707e+17, 1.297991118534771e+17, 1.297991118575395e+17, 1.297991118616019e+17, 1.297991118655082e+17, 1.297991118695707e+17, 1.297991118736333e+17, 1.297991118775395e+17, 1.29799111881602e+17, 1.297991118856645e+17, 1.297991118895708e+17, 1.297991118936333e+17, 1.297991118976957e+17, 1.297991119017582e+17, 1.297991119056645e+17, 1.29799111909727e+17, 1.297991119137896e+17, 1.297991119176957e+17, 1.297991119217582e+17, 1.297991119258208e+17, 1.297991119298833e+17, 1.297991119337894e+17, 1.29799111937852e+17, 1.297991119419145e+17, 1.297991119458208e+17, 1.297991119498833e+17, 1.297991119539457e+17, 1.29799111957852e+17, 1.297991119619145e+17, 1.29799111965977e+17, 1.297991119700396e+17, 1.297991119739457e+17, 1.297991119780083e+17, 1.297991119820708e+17, 1.297991119859771e+17, 1.297991119900394e+17, 1.29799111994102e+17, 1.297991119981645e+17, 1.297991120020707e+17, 1.297991120061332e+17, 1.297991120101958e+17, 1.29799112014102e+17, 1.297991120181646e+17, 1.297991120222269e+17, 1.297991120261332e+17, 1.297991120301958e+17, 1.297991120342582e+17, 1.297991120383208e+17, 1.297991120422269e+17, 1.297991120462895e+17, 1.29799112050352e+17, 1.297991120542583e+17, 1.297991120583208e+17, 1.297991120623832e+17, 1.297991120662895e+17, 1.29799112070352e+17, 1.297991120744145e+17, 1.297991120783208e+17, 1.297991120823832e+17, 1.297991120864457e+17, 1.297991120905083e+17, 1.297991120944145e+17, 1.297991120984769e+17, 1.297991121025395e+17, 1.297991121064457e+17, 1.297991121105083e+17, 1.297991121145708e+17, 1.297991121186332e+17, 1.297991121225395e+17, 1.29799112126602e+17, 1.297991121306644e+17, 1.297991121345708e+17, 1.297991121386332e+17, 1.297991121426958e+17, 1.29799112146602e+17, 1.297991121506646e+17, 1.29799112154727e+17, 1.297991121587895e+17, 1.297991121626958e+17, 1.297991121667581e+17, 1.297991121708207e+17, 1.29799112174727e+17, 1.297991121787895e+17, 1.297991121828521e+17, 1.297991121869146e+17, 1.297991121908207e+17, 1.297991121948833e+17, 1.297991121989457e+17, 1.29799112202852e+17, 1.297991122069144e+17, 1.29799112210977e+17, 1.297991122148833e+17, 1.297991122189458e+17, 1.297991122230083e+17, 1.297991122270707e+17, 1.29799112230977e+17, 1.297991122350395e+17, 1.29799112239102e+17, 1.297991122430083e+17, 1.297991122470707e+17, 1.297991122511332e+17, 1.297991122550396e+17, 1.29799112259102e+17, 1.297991122631645e+17, 1.297991122670707e+17, 1.297991122711332e+17, 1.297991122751958e+17, 1.297991122792582e+17, 1.297991122831645e+17, 1.29799112287227e+17, 1.297991122912895e+17, 1.297991122951958e+17, 1.297991122992582e+17, 1.297991123033207e+17, 1.297991123073833e+17, 1.297991123112895e+17, 1.297991123153521e+17, 1.297991123194145e+17, 1.297991123233207e+17, 1.297991123273833e+17, 1.297991123314458e+17, 1.297991123353521e+17, 1.297991123394145e+17, 1.29799112343477e+17, 1.297991123475396e+17, 1.297991123514458e+17, 1.297991123555082e+17, 1.297991123595708e+17, 1.29799112363477e+17, 1.297991123675395e+17, 1.29799112371602e+17, 1.297991123756645e+17, 1.297991123795708e+17, 1.297991123836333e+17, 1.297991123876957e+17, 1.297991123916019e+17, 1.297991123956645e+17, 1.29799112399727e+17, 1.297991124036332e+17, 1.297991124076957e+17, 1.297991124117583e+17, 1.297991124158207e+17, 1.297991124197271e+17, 1.297991124237894e+17, 1.29799112427852e+17, 1.297991124317583e+17, 1.297991124358207e+17, 1.297991124398833e+17, 1.297991124437894e+17, 1.29799112447852e+17, 1.297991124519145e+17, 1.297991124558208e+17, 1.297991124598833e+17, 1.297991124639457e+17, 1.297991124680082e+17, 1.297991124719145e+17, 1.29799112475977e+17, 1.297991124800396e+17, 1.297991124839457e+17, 1.297991124880082e+17, 1.297991124920708e+17, 1.297991124961332e+17, 1.297991125000396e+17, 1.29799112504102e+17, 1.297991125081645e+17, 1.297991125120708e+17, 1.297991125161332e+17, 1.297991125201957e+17, 1.29799112524102e+17, 1.297991125281645e+17, 1.297991125322269e+17, 1.297991125362895e+17, 1.297991125401957e+17, 1.297991125442583e+17, 1.297991125483208e+17, 1.297991125522271e+17, 1.297991125562895e+17, 1.29799112560352e+17, 1.297991125644145e+17, 1.297991125683206e+17, 1.297991125723832e+17, 1.297991125764458e+17, 1.29799112580352e+17, 1.297991125844146e+17, 1.297991125884771e+17, 1.297991125923832e+17, 1.297991125964458e+17, 1.297991126005082e+17, 1.297991126045708e+17, 1.297991126084769e+17, 1.297991126125395e+17, 1.29799112616602e+17, 1.297991126205083e+17, 1.297991126245708e+17, 1.297991126286333e+17, 1.297991126325395e+17, 1.29799112636602e+17, 1.297991126406644e+17, 1.297991126445708e+17, 1.297991126486332e+17, 1.297991126526957e+17, 1.297991126567583e+17, 1.297991126606644e+17, 1.29799112664727e+17, 1.297991126687895e+17, 1.297991126726957e+17, 1.297991126767583e+17, 1.297991126808207e+17, 1.297991126848832e+17, 1.297991126887895e+17, 1.29799112692852e+17, 1.297991126969144e+17, 1.297991127008207e+17, 1.297991127048832e+17, 1.297991127089458e+17, 1.29799112712852e+17, 1.297991127169146e+17, 1.29799112720977e+17, 1.297991127250395e+17, 1.297991127289458e+17, 1.297991127330083e+17, 1.297991127370707e+17, 1.29799112740977e+17, 1.297991127450395e+17, 1.297991127491021e+17, 1.297991127531645e+17, 1.297991127570707e+17, 1.297991127611333e+17, 1.297991127651958e+17, 1.29799112769102e+17, 1.297991127731645e+17, 1.29799112777227e+17, 1.297991127811333e+17, 1.297991127851958e+17, 1.297991127892582e+17, 1.297991127933208e+17, 1.29799112797227e+17, 1.297991128012895e+17, 1.297991128053521e+17, 1.297991128092582e+17, 1.297991128133208e+17, 1.297991128173832e+17, 1.297991128212896e+17, 1.297991128253519e+17, 1.297991128294145e+17, 1.297991128333208e+17, 1.297991128373832e+17, 1.297991128414458e+17, 1.297991128455084e+17, 1.297991128494145e+17, 1.29799112853477e+17, 1.297991128575395e+17, 1.297991128614458e+17, 1.297991128655082e+17, 1.297991128695707e+17, 1.297991128736333e+17, 1.297991128775395e+17, 1.29799112881602e+17, 1.297991128856645e+17, 1.297991128895707e+17, 1.297991128936333e+17, 1.297991128976957e+17, 1.29799112901602e+17, 1.297991129056645e+17, 1.29799112909727e+17, 1.297991129137896e+17, 1.297991129176957e+17, 1.297991129217582e+17, 1.297991129258208e+17, 1.29799112929727e+17, 1.297991129337894e+17, 1.29799112937852e+17, 1.297991129419145e+17, 1.297991129458208e+17, 1.297991129498833e+17, 1.297991129539457e+17, 1.29799112957852e+17, 1.297991129619145e+17, 1.29799112965977e+17, 1.297991129698831e+17, 1.297991129739457e+17, 1.297991129780083e+17, 1.297991129820707e+17, 1.297991129859771e+17, 1.297991129900396e+17, 1.29799112994102e+17, 1.297991129980083e+17, 1.297991130020707e+17, 1.297991130061332e+17, 1.297991130100394e+17, 1.29799113014102e+17, 1.297991130181645e+17, 1.297991130220708e+17, 1.297991130261332e+17, 1.297991130301958e+17, 1.297991130342582e+17, 1.297991130381645e+17, 1.297991130422269e+17, 1.297991130462895e+17, 1.297991130501957e+17, 1.297991130542582e+17, 1.297991130583208e+17, 1.297991130623832e+17, 1.297991130662895e+17, 1.29799113070352e+17, 1.297991130744145e+17, 1.297991130783208e+17, 1.297991130823832e+17, 1.297991130864457e+17, 1.29799113090352e+17, 1.297991130944145e+17, 1.297991130984769e+17, 1.297991131025395e+17, 1.297991131064457e+17, 1.297991131105083e+17, 1.297991131145708e+17, 1.297991131184771e+17, 1.297991131225395e+17, 1.29799113126602e+17, 1.297991131306644e+17, 1.297991131345708e+17, 1.297991131386332e+17, 1.297991131426958e+17, 1.29799113146602e+17, 1.297991131506646e+17, 1.29799113154727e+17, 1.297991131586332e+17, 1.297991131626958e+17, 1.297991131667583e+17, 1.297991131708207e+17, 1.29799113174727e+17, 1.297991131787895e+17, 1.29799113182852e+17, 1.297991131867583e+17, 1.297991131908207e+17, 1.297991131948833e+17, 1.297991131987895e+17, 1.29799113202852e+17, 1.297991132069146e+17, 1.297991132108207e+17, 1.297991132148833e+17, 1.297991132189457e+17, 1.297991132230083e+17, 1.297991132269144e+17, 1.29799113230977e+17, 1.297991132350395e+17, 1.297991132389457e+17, 1.297991132430083e+17, 1.297991132470708e+17, 1.297991132511332e+17, 1.297991132550395e+17, 1.29799113259102e+17, 1.297991132631644e+17, 1.297991132670707e+17, 1.297991132711332e+17, 1.297991132751958e+17, 1.29799113279102e+17, 1.297991132831645e+17, 1.29799113287227e+17, 1.297991132912895e+17, 1.297991132951958e+17, 1.297991132992582e+17, 1.297991133033207e+17, 1.29799113307227e+17, 1.297991133112895e+17, 1.297991133153521e+17, 1.297991133194145e+17, 1.297991133233207e+17, 1.297991133273833e+17, 1.297991133314458e+17, 1.297991133353519e+17, 1.297991133394145e+17, 1.29799113343477e+17, 1.297991133473833e+17, 1.297991133514458e+17, 1.297991133555082e+17, 1.297991133595708e+17, 1.29799113363477e+17, 1.297991133675395e+17, 1.29799113371602e+17, 1.297991133755082e+17, 1.297991133795708e+17, 1.297991133836332e+17, 1.297991133875396e+17, 1.29799113391602e+17, 1.297991133956645e+17, 1.297991133995708e+17, 1.297991134036332e+17, 1.297991134076957e+17, 1.297991134117583e+17, 1.297991134156645e+17, 1.29799113419727e+17, 1.297991134237896e+17, 1.297991134276957e+17, 1.297991134317583e+17, 1.297991134358207e+17, 1.297991134398833e+17, 1.297991134437894e+17, 1.29799113447852e+17, 1.297991134519145e+17, 1.297991134558208e+17, 1.297991134598833e+17, 1.297991134639457e+17, 1.29799113467852e+17, 1.297991134719145e+17, 1.29799113475977e+17, 1.297991134800396e+17, 1.297991134839457e+17, 1.297991134880082e+17, 1.297991134920708e+17, 1.29799113495977e+17, 1.297991135000394e+17, 1.29799113504102e+17, 1.297991135081645e+17, 1.297991135120708e+17, 1.297991135161332e+17, 1.297991135201957e+17, 1.29799113524102e+17, 1.297991135281645e+17, 1.297991135322269e+17, 1.297991135361332e+17, 1.297991135401957e+17, 1.297991135442583e+17, 1.297991135483208e+17, 1.297991135522271e+17, 1.297991135562895e+17, 1.29799113560352e+17, 1.297991135642583e+17, 1.297991135683208e+17, 1.297991135723832e+17, 1.297991135762895e+17, 1.29799113580352e+17, 1.297991135844145e+17, 1.297991135883208e+17, 1.297991135923832e+17, 1.297991135964458e+17, 1.297991136005082e+17, 1.297991136044145e+17, 1.297991136084771e+17, 1.297991136125395e+17, 1.297991136164458e+17, 1.297991136205083e+17, 1.297991136245708e+17, 1.297991136286332e+17, 1.297991136325395e+17, 1.29799113636602e+17, 1.297991136406644e+17, 1.297991136445708e+17, 1.297991136486333e+17, 1.297991136526957e+17, 1.297991136566021e+17, 1.297991136606644e+17, 1.297991136647269e+17, 1.297991136687895e+17, 1.297991136726957e+17, 1.297991136767583e+17, 1.297991136808209e+17, 1.29799113684727e+17, 1.297991136887895e+17, 1.29799113692852e+17, 1.297991136969144e+17, 1.297991137008207e+17, 1.297991137048832e+17, 1.297991137089458e+17, 1.29799113712852e+17, 1.297991137169146e+17, 1.29799113720977e+17, 1.297991137248832e+17, 1.297991137289458e+17, 1.297991137330083e+17, 1.297991137370707e+17, 1.29799113740977e+17, 1.297991137450395e+17, 1.297991137491021e+17, 1.297991137530083e+17, 1.297991137570707e+17, 1.297991137611333e+17, 1.297991137650395e+17, 1.29799113769102e+17, 1.297991137731645e+17, 1.297991137770707e+17, 1.297991137811333e+17, 1.297991137851958e+17, 1.297991137892582e+17, 1.297991137931645e+17, 1.29799113797227e+17, 1.297991138012895e+17, 1.297991138051956e+17, 1.297991138092582e+17, 1.297991138133208e+17, 1.297991138173832e+17, 1.297991138212896e+17, 1.297991138253521e+17, 1.297991138294144e+17, 1.297991138333208e+17, 1.297991138373832e+17, 1.297991138414458e+17, 1.297991138453519e+17, 1.297991138494145e+17, 1.29799113853477e+17, 1.297991138575395e+17, 1.297991138614458e+17, 1.297991138655082e+17, 1.297991138695707e+17, 1.29799113873477e+17, 1.297991138775395e+17, 1.29799113881602e+17, 1.297991138856645e+17, 1.297991138895707e+17, 1.297991138936333e+17, 1.297991138976957e+17, 1.297991139016019e+17, 1.297991139056645e+17, 1.29799113909727e+17, 1.297991139136333e+17, 1.297991139176957e+17, 1.297991139217582e+17, 1.297991139258208e+17, 1.29799113929727e+17, 1.297991139337894e+17, 1.29799113937852e+17, 1.297991139417582e+17, 1.297991139458208e+17, 1.297991139498833e+17, 1.297991139537896e+17, 1.29799113957852e+17, 1.297991139619145e+17, 1.297991139658208e+17, 1.297991139698833e+17, 1.297991139739457e+17, 1.297991139780083e+17, 1.297991139819145e+17, 1.297991139859771e+17, 1.297991139900396e+17, 1.297991139939457e+17, 1.297991139980083e+17, 1.297991140020707e+17, 1.297991140061332e+17, 1.297991140100396e+17, 1.29799114014102e+17, 1.297991140181645e+17, 1.297991140220708e+17, 1.297991140261332e+17, 1.297991140301957e+17, 1.29799114034102e+17, 1.297991140381645e+17, 1.297991140422269e+17, 1.297991140462895e+17, 1.297991140501958e+17, 1.297991140542582e+17, 1.297991140583208e+17, 1.297991140622269e+17, 1.297991140662894e+17, 1.29799114070352e+17, 1.297991140744145e+17, 1.297991140783208e+17, 1.297991140823834e+17, 1.297991140864457e+17, 1.29799114090352e+17, 1.297991140944145e+17, 1.297991140984769e+17, 1.297991141023832e+17, 1.297991141064457e+17, 1.297991141105083e+17, 1.297991141145708e+17, 1.297991141184771e+17, 1.297991141225395e+17, 1.29799114126602e+17, 1.297991141305083e+17, 1.297991141345708e+17, 1.297991141386332e+17, 1.297991141425395e+17, 1.29799114146602e+17, 1.297991141506646e+17, 1.297991141545708e+17, 1.297991141586332e+17, 1.297991141626958e+17, 1.297991141667583e+17, 1.297991141706644e+17, 1.29799114174727e+17, 1.297991141787895e+17, 1.297991141826958e+17, 1.297991141867583e+17, 1.297991141908207e+17, 1.297991141948832e+17, 1.297991141987895e+17, 1.29799114202852e+17, 1.297991142069146e+17, 1.297991142108207e+17, 1.297991142148833e+17, 1.297991142189457e+17, 1.297991142228521e+17, 1.297991142269146e+17, 1.297991142309769e+17, 1.297991142350395e+17, 1.297991142389457e+17, 1.297991142430083e+17, 1.297991142470708e+17, 1.29799114250977e+17, 1.297991142550395e+17, 1.29799114259102e+17, 1.297991142631644e+17, 1.297991142670708e+17, 1.297991142711332e+17, 1.297991142751958e+17, 1.29799114279102e+17, 1.297991142831645e+17, 1.29799114287227e+17, 1.297991142911332e+17, 1.297991142951958e+17, 1.297991142992582e+17, 1.297991143033207e+17, 1.29799114307227e+17, 1.297991143112895e+17, 1.297991143153521e+17, 1.297991143192582e+17, 1.297991143233207e+17, 1.297991143273833e+17, 1.297991143312895e+17, 1.297991143353519e+17, 1.297991143394145e+17, 1.297991143433207e+17, 1.297991143473833e+17, 1.297991143514458e+17, 1.297991143555082e+17, 1.297991143594145e+17, 1.29799114363477e+17, 1.297991143675395e+17, 1.297991143714458e+17, 1.297991143755082e+17, 1.297991143795708e+17, 1.297991143836333e+17, 1.297991143875396e+17, 1.29799114391602e+17, 1.297991143956644e+17, 1.297991143995708e+17, 1.297991144036332e+17, 1.297991144076957e+17, 1.29799114411602e+17, 1.297991144156645e+17, 1.29799114419727e+17, 1.297991144237896e+17, 1.297991144276957e+17, 1.297991144317583e+17, 1.297991144358207e+17, 1.29799114439727e+17, 1.297991144437896e+17, 1.29799114447852e+17, 1.297991144519145e+17, 1.297991144558207e+17, 1.297991144598833e+17, 1.297991144639457e+17, 1.29799114467852e+17, 1.297991144719145e+17, 1.29799114475977e+17, 1.297991144798833e+17, 1.297991144839459e+17, 1.297991144880082e+17, 1.297991144920708e+17, 1.29799114495977e+17, 1.297991145000394e+17, 1.29799114504102e+17, 1.297991145080082e+17, 1.297991145120708e+17, 1.297991145161332e+17, 1.297991145200396e+17, 1.29799114524102e+17, 1.297991145281645e+17, 1.297991145320708e+17, 1.297991145361332e+17, 1.297991145401957e+17, 1.297991145442583e+17, 1.297991145481645e+17, 1.297991145522271e+17, 1.297991145562895e+17, 1.297991145601957e+17, 1.297991145642583e+17, 1.297991145683208e+17, 1.297991145723832e+17, 1.297991145762895e+17, 1.29799114580352e+17, 1.297991145844145e+17, 1.297991145883208e+17, 1.297991145923832e+17, 1.297991145964458e+17, 1.29799114600352e+17, 1.297991146044145e+17, 1.297991146084771e+17, 1.297991146125395e+17, 1.297991146164458e+17, 1.297991146205082e+17, 1.297991146245708e+17, 1.297991146284771e+17, 1.297991146325395e+17, 1.29799114636602e+17, 1.297991146406646e+17, 1.297991146445708e+17, 1.297991146486333e+17, 1.297991146526957e+17, 1.29799114656602e+17, 1.297991146606644e+17, 1.297991146647269e+17, 1.297991146686333e+17, 1.297991146726957e+17, 1.297991146767583e+17, 1.297991146808209e+17, 1.29799114684727e+17, 1.297991146887895e+17, 1.29799114692852e+17, 1.297991146967583e+17, 1.297991147008207e+17, 1.297991147048832e+17, 1.297991147087895e+17, 1.29799114712852e+17, 1.297991147169146e+17, 1.297991147208207e+17, 1.297991147248832e+17, 1.297991147289458e+17, 1.297991147330083e+17, 1.297991147369144e+17, 1.29799114740977e+17, 1.297991147450395e+17, 1.297991147489458e+17, 1.297991147530083e+17, 1.297991147570707e+17, 1.297991147611333e+17, 1.297991147650395e+17, 1.29799114769102e+17, 1.297991147731645e+17, 1.297991147770707e+17, 1.297991147811333e+17, 1.297991147851958e+17, 1.297991147891021e+17, 1.297991147931645e+17, 1.29799114797227e+17, 1.297991148012895e+17, 1.297991148051956e+17, 1.297991148092582e+17, 1.297991148133208e+17, 1.29799114817227e+17, 1.297991148212895e+17, 1.297991148253521e+17, 1.297991148294144e+17, 1.297991148333208e+17, 1.297991148373832e+17, 1.297991148414458e+17, 1.297991148453521e+17, 1.297991148494145e+17, 1.29799114853477e+17, 1.297991148573832e+17, 1.297991148614458e+17, 1.297991148655082e+17, 1.297991148695707e+17, 1.29799114873477e+17, 1.297991148775395e+17, 1.29799114881602e+17, 1.297991148855084e+17, 1.297991148895707e+17, 1.297991148936333e+17, 1.297991148975395e+17, 1.297991149016019e+17, 1.297991149056645e+17, 1.297991149095707e+17, 1.297991149136333e+17, 1.297991149176957e+17, 1.297991149217582e+17, 1.297991149256645e+17, 1.29799114929727e+17, 1.297991149337894e+17, 1.297991149376957e+17, 1.297991149417582e+17, 1.297991149458208e+17, 1.297991149498833e+17, 1.297991149537896e+17, 1.29799114957852e+17, 1.297991149619145e+17, 1.297991149658208e+17, 1.297991149698833e+17, 1.297991149739457e+17, 1.29799114977852e+17, 1.297991149819145e+17, 1.29799114985977e+17, 1.297991149900396e+17, 1.297991149939457e+17, 1.297991149980083e+17, 1.297991150020708e+17, 1.29799115005977e+17, 1.297991150100396e+17, 1.29799115014102e+17, 1.297991150181645e+17, 1.297991150220707e+17, 1.297991150261332e+17, 1.297991150301957e+17, 1.29799115034102e+17, 1.297991150381645e+17, 1.297991150422271e+17, 1.297991150461332e+17, 1.297991150501958e+17, 1.297991150542582e+17, 1.297991150583208e+17, 1.297991150622269e+17, 1.297991150662894e+17, 1.29799115070352e+17, 1.297991150742582e+17, 1.297991150783208e+17, 1.297991150823834e+17, 1.297991150862895e+17, 1.29799115090352e+17, 1.297991150944145e+17, 1.297991150983208e+17, 1.297991151023832e+17, 1.297991151064457e+17, 1.297991151105083e+17, 1.297991151144145e+17, 1.297991151184771e+17, 1.297991151225395e+17, 1.297991151264457e+17, 1.297991151305083e+17, 1.297991151345708e+17, 1.297991151386332e+17, 1.297991151425395e+17, 1.29799115146602e+17, 1.297991151506644e+17, 1.297991151545708e+17, 1.297991151586332e+17, 1.297991151626958e+17, 1.29799115166602e+17, 1.297991151706644e+17, 1.29799115174727e+17, 1.297991151787895e+17, 1.297991151826958e+17, 1.297991151867583e+17, 1.297991151908207e+17, 1.29799115194727e+17, 1.297991151987895e+17, 1.29799115202852e+17, 1.297991152069146e+17, 1.297991152108207e+17, 1.297991152148833e+17, 1.297991152189458e+17, 1.29799115222852e+17, 1.297991152269146e+17, 1.297991152309769e+17, 1.297991152348833e+17, 1.297991152389457e+17, 1.297991152430083e+17, 1.297991152470708e+17, 1.29799115250977e+17, 1.297991152550395e+17, 1.297991152591021e+17, 1.297991152630083e+17, 1.297991152670707e+17, 1.297991152711332e+17, 1.297991152750395e+17, 1.29799115279102e+17, 1.297991152831645e+17, 1.297991152870708e+17, 1.297991152911332e+17, 1.297991152951958e+17, 1.297991152992582e+17, 1.297991153031644e+17, 1.29799115307227e+17, 1.297991153112895e+17, 1.297991153151958e+17, 1.297991153192582e+17, 1.297991153233207e+17, 1.297991153273833e+17, 1.297991153312895e+17, 1.297991153353519e+17, 1.297991153394145e+17, 1.297991153433207e+17, 1.297991153473833e+17, 1.297991153514458e+17, 1.297991153553521e+17, 1.297991153594145e+17, 1.29799115363477e+17, 1.297991153675395e+17, 1.297991153714458e+17, 1.297991153755082e+17, 1.297991153795708e+17, 1.29799115383477e+17, 1.297991153875395e+17, 1.29799115391602e+17, 1.297991153956644e+17, 1.297991153995708e+17, 1.297991154036333e+17, 1.297991154076957e+17, 1.29799115411602e+17, 1.297991154156645e+17, 1.29799115419727e+17, 1.297991154236332e+17, 1.297991154276957e+17, 1.297991154317582e+17, 1.297991154358207e+17, 1.29799115439727e+17, 1.297991154437896e+17, 1.29799115447852e+17, 1.297991154517583e+17, 1.297991154558207e+17, 1.297991154598833e+17, 1.297991154637896e+17, 1.297991154678519e+17, 1.297991154719145e+17, 1.297991154758207e+17, 1.297991154798833e+17, 1.297991154839459e+17, 1.297991154880082e+17, 1.297991154919145e+17, 1.29799115495977e+17, 1.297991155000394e+17, 1.297991155039457e+17, 1.297991155080082e+17, 1.297991155120708e+17, 1.297991155161332e+17, 1.297991155200396e+17, 1.29799115524102e+17, 1.297991155281645e+17, 1.297991155320708e+17, 1.297991155361332e+17, 1.297991155401957e+17, 1.29799115544102e+17, 1.297991155481645e+17, 1.297991155522269e+17, 1.297991155562895e+17, 1.297991155601957e+17, 1.297991155642583e+17, 1.297991155683208e+17, 1.297991155722269e+17, 1.297991155762895e+17, 1.29799115580352e+17, 1.297991155844145e+17, 1.297991155883208e+17, 1.297991155923832e+17, 1.297991155964457e+17, 1.29799115600352e+17, 1.297991156044145e+17, 1.297991156084771e+17, 1.297991156123832e+17, 1.297991156164458e+17, 1.297991156205083e+17, 1.297991156245708e+17, 1.297991156284771e+17, 1.297991156325394e+17, 1.29799115636602e+17, 1.297991156405082e+17, 1.297991156445708e+17, 1.297991156486333e+17, 1.297991156525395e+17, 1.29799115656602e+17, 1.297991156606646e+17, 1.297991156645708e+17, 1.297991156686332e+17, 1.297991156726957e+17, 1.297991156767583e+17, 1.297991156806644e+17, 1.29799115684727e+17, 1.297991156887895e+17, 1.297991156926957e+17, 1.297991156967583e+17, 1.297991157008207e+17, 1.297991157048832e+17, 1.297991157087895e+17, 1.29799115712852e+17, 1.297991157169144e+17, 1.297991157208207e+17, 1.297991157248832e+17, 1.297991157289458e+17, 1.29799115732852e+17, 1.297991157369144e+17, 1.29799115740977e+17, 1.297991157450395e+17, 1.297991157489458e+17, 1.297991157530083e+17, 1.297991157570707e+17, 1.29799115760977e+17, 1.297991157650395e+17, 1.29799115769102e+17, 1.297991157731645e+17, 1.297991157770707e+17, 1.297991157811333e+17, 1.297991157851958e+17, 1.297991157891021e+17, 1.297991157931645e+17, 1.297991157972269e+17, 1.297991158011333e+17, 1.297991158051958e+17, 1.297991158092582e+17, 1.297991158133208e+17, 1.29799115817227e+17, 1.297991158212895e+17, 1.297991158253521e+17, 1.297991158292582e+17, 1.297991158333207e+17, 1.297991158373833e+17, 1.297991158412895e+17, 1.297991158453521e+17, 1.297991158494145e+17, 1.297991158533208e+17, 1.297991158573832e+17, 1.297991158614458e+17, 1.297991158655082e+17, 1.297991158694144e+17, 1.29799115873477e+17, 1.297991158775396e+17, 1.297991158814458e+17, 1.297991158855084e+17, 1.297991158895707e+17, 1.297991158936333e+17, 1.297991158975395e+17, 1.297991159016019e+17, 1.297991159056645e+17, 1.297991159095707e+17, 1.297991159136333e+17, 1.297991159176959e+17, 1.29799115921602e+17, 1.297991159256645e+17, 1.29799115929727e+17, 1.297991159337894e+17, 1.297991159376957e+17, 1.297991159417582e+17, 1.297991159458208e+17, 1.29799115949727e+17, 1.297991159537896e+17, 1.29799115957852e+17, 1.297991159619145e+17, 1.297991159658208e+17, 1.297991159698833e+17, 1.297991159739457e+17, 1.29799115977852e+17, 1.297991159819145e+17, 1.29799115985977e+17, 1.297991159898833e+17, 1.297991159939457e+17, 1.297991159980082e+17, 1.297991160020708e+17, 1.29799116005977e+17, 1.297991160100396e+17, 1.29799116014102e+17, 1.297991160180083e+17, 1.297991160220708e+17, 1.297991160261332e+17, 1.297991160300396e+17, 1.297991160341019e+17, 1.297991160381645e+17, 1.297991160420707e+17, 1.297991160461332e+17, 1.297991160501958e+17, 1.297991160542582e+17, 1.297991160581645e+17, 1.297991160622271e+17, 1.297991160662894e+17, 1.297991160701957e+17, 1.297991160742582e+17, 1.297991160783208e+17, 1.297991160823834e+17, 1.297991160862895e+17, 1.29799116090352e+17, 1.297991160944146e+17, 1.297991160983208e+17, 1.297991161023832e+17, 1.297991161064457e+17, 1.29799116110352e+17, 1.297991161144145e+17, 1.297991161184771e+17, 1.297991161225395e+17, 1.297991161264457e+17, 1.297991161305083e+17, 1.297991161345708e+17, 1.297991161384769e+17, 1.297991161425395e+17, 1.29799116146602e+17, 1.297991161506644e+17, 1.297991161545708e+17, 1.297991161586332e+17, 1.297991161626957e+17, 1.29799116166602e+17, 1.297991161706644e+17, 1.29799116174727e+17, 1.297991161786332e+17, 1.297991161826958e+17, 1.297991161867583e+17, 1.297991161908207e+17, 1.29799116194727e+17, 1.297991161987895e+17, 1.29799116202852e+17, 1.297991162067583e+17, 1.297991162108207e+17, 1.297991162148833e+17, 1.297991162187895e+17, 1.29799116222852e+17, 1.297991162269146e+17, 1.297991162308207e+17, 1.297991162348832e+17, 1.297991162389458e+17, 1.297991162430083e+17, 1.297991162469146e+17, 1.29799116250977e+17, 1.297991162550395e+17, 1.297991162589457e+17, 1.297991162630083e+17, 1.297991162670707e+17, 1.297991162711332e+17, 1.297991162750395e+17, 1.297991162791021e+17, 1.297991162831645e+17, 1.297991162870708e+17, 1.297991162911332e+17, 1.297991162951958e+17, 1.29799116299102e+17, 1.297991163031644e+17, 1.29799116307227e+17, 1.297991163112895e+17, 1.297991163151958e+17, 1.297991163192584e+17, 1.297991163233207e+17, 1.29799116327227e+17, 1.297991163312895e+17, 1.297991163353519e+17, 1.297991163394145e+17, 1.297991163433207e+17, 1.297991163473833e+17, 1.297991163514458e+17, 1.297991163553521e+17, 1.297991163594145e+17, 1.29799116363477e+17, 1.297991163673833e+17, 1.297991163714458e+17, 1.297991163755082e+17, 1.297991163795708e+17, 1.29799116383477e+17, 1.297991163875395e+17, 1.29799116391602e+17, 1.297991163955082e+17, 1.297991163995707e+17, 1.297991164036333e+17, 1.297991164075395e+17, 1.29799116411602e+17, 1.297991164156645e+17, 1.297991164195708e+17, 1.297991164236333e+17, 1.297991164276957e+17, 1.297991164317582e+17, 1.297991164356645e+17, 1.29799116439727e+17, 1.297991164437896e+17, 1.297991164476957e+17, 1.297991164517583e+17, 1.297991164558207e+17, 1.297991164598833e+17, 1.297991164637896e+17, 1.297991164678519e+17, 1.297991164719145e+17, 1.297991164758207e+17, 1.297991164798833e+17, 1.297991164839459e+17, 1.29799116487852e+17, 1.297991164919145e+17, 1.297991164959771e+17, 1.297991165000394e+17, 1.297991165039457e+17, 1.297991165080082e+17, 1.297991165120708e+17, 1.29799116515977e+17, 1.297991165200396e+17, 1.29799116524102e+17, 1.297991165281645e+17, 1.297991165320708e+17, 1.297991165361332e+17, 1.297991165401957e+17, 1.29799116544102e+17, 1.297991165481645e+17, 1.297991165522269e+17, 1.297991165561332e+17, 1.297991165601957e+17, 1.297991165642583e+17, 1.297991165683208e+17, 1.297991165722269e+17, 1.297991165762895e+17, 1.29799116580352e+17, 1.297991165842583e+17, 1.297991165883208e+17, 1.297991165923832e+17, 1.297991165962895e+17, 1.29799116600352e+17, 1.297991166044145e+17, 1.297991166083208e+17, 1.297991166123832e+17, 1.297991166164458e+17, 1.297991166205083e+17, 1.297991166244145e+17, 1.297991166284771e+17, 1.297991166325394e+17, 1.297991166364458e+17, 1.297991166405083e+17, 1.297991166445708e+17, 1.297991166486333e+17, 1.297991166525395e+17, 1.29799116656602e+17, 1.297991166606646e+17, 1.297991166645708e+17, 1.297991166686332e+17, 1.297991166726957e+17, 1.29799116676602e+17, 1.297991166806646e+17, 1.29799116684727e+17, 1.297991166887895e+17, 1.297991166926957e+17, 1.297991166967583e+17, 1.297991167008207e+17, 1.297991167047269e+17, 1.297991167087895e+17, 1.29799116712852e+17, 1.297991167169144e+17, 1.297991167208209e+17, 1.297991167248832e+17, 1.297991167289458e+17, 1.29799116732852e+17, 1.297991167369144e+17, 1.29799116740977e+17, 1.297991167448832e+17, 1.297991167489458e+17, 1.297991167530083e+17, 1.297991167570707e+17, 1.29799116760977e+17, 1.297991167650395e+17, 1.29799116769102e+17, 1.297991167730083e+17, 1.297991167770707e+17, 1.297991167811333e+17, 1.297991167850395e+17, 1.29799116789102e+17, 1.297991167931645e+17, 1.297991167970707e+17, 1.297991168011333e+17, 1.297991168051958e+17, 1.297991168092582e+17, 1.297991168131645e+17, 1.29799116817227e+17, 1.297991168212895e+17, 1.297991168251958e+17, 1.297991168292582e+17, 1.297991168333207e+17, 1.297991168373833e+17, 1.297991168412895e+17, 1.297991168453521e+17, 1.297991168494145e+17, 1.297991168533208e+17, 1.297991168573833e+17, 1.297991168614458e+17, 1.297991168653521e+17, 1.297991168694144e+17, 1.29799116873477e+17, 1.297991168775396e+17, 1.297991168814458e+17, 1.297991168855084e+17, 1.297991168895707e+17, 1.29799116893477e+17, 1.297991168975396e+17, 1.297991169016019e+17, 1.297991169056645e+17, 1.297991169095707e+17, 1.297991169136333e+17, 1.297991169176957e+17, 1.29799116921602e+17, 1.297991169256645e+17, 1.29799116929727e+17, 1.297991169336333e+17, 1.297991169376957e+17, 1.297991169417582e+17, 1.297991169458208e+17, 1.29799116949727e+17, 1.297991169537894e+17, 1.29799116957852e+17, 1.297991169617582e+17, 1.297991169658208e+17, 1.297991169698833e+17, 1.297991169737894e+17, 1.29799116977852e+17, 1.297991169819145e+17, 1.297991169858208e+17, 1.297991169898833e+17, 1.297991169939457e+17, 1.297991169980082e+17, 1.297991170019145e+17, 1.29799117005977e+17, 1.297991170100396e+17, 1.297991170139457e+17, 1.297991170180083e+17, 1.297991170220708e+17, 1.297991170261332e+17, 1.297991170300396e+17, 1.297991170341019e+17, 1.297991170381645e+17, 1.297991170420708e+17, 1.297991170461332e+17, 1.297991170501958e+17, 1.29799117054102e+17, 1.297991170581645e+17, 1.297991170622271e+17, 1.297991170662894e+17, 1.297991170701957e+17, 1.297991170742582e+17, 1.297991170783208e+17, 1.297991170822271e+17, 1.297991170862895e+17, 1.29799117090352e+17, 1.297991170944146e+17, 1.297991170983208e+17, 1.297991171023832e+17, 1.297991171064457e+17, 1.29799117110352e+17, 1.297991171144146e+17, 1.297991171184769e+17, 1.297991171223834e+17, 1.297991171264457e+17, 1.297991171305083e+17, 1.297991171345708e+17, 1.297991171384769e+17, 1.297991171425395e+17, 1.29799117146602e+17, 1.297991171505083e+17, 1.297991171545708e+17, 1.297991171586332e+17, 1.297991171625395e+17, 1.29799117166602e+17, 1.297991171706644e+17, 1.297991171745708e+17, 1.297991171786332e+17, 1.297991171826958e+17, 1.297991171867583e+17, 1.297991171906644e+17, 1.29799117194727e+17, 1.297991171987895e+17, 1.297991172026958e+17, 1.297991172067583e+17, 1.297991172108207e+17, 1.297991172148833e+17, 1.297991172187895e+17, 1.29799117222852e+17, 1.297991172269146e+17, 1.297991172308207e+17, 1.297991172348832e+17, 1.297991172389458e+17, 1.29799117242852e+17, 1.297991172469146e+17, 1.29799117250977e+17, 1.297991172550395e+17, 1.297991172589458e+17, 1.297991172630083e+17, 1.297991172670707e+17, 1.297991172709769e+17, 1.297991172750395e+17, 1.297991172791021e+17, 1.297991172831644e+17, 1.297991172870708e+17, 1.297991172911332e+17, 1.297991172951958e+17, 1.297991172991021e+17, 1.297991173031644e+17, 1.29799117307227e+17, 1.297991173111332e+17, 1.297991173151958e+17, 1.297991173192582e+17, 1.297991173233207e+17, 1.29799117327227e+17, 1.297991173312895e+17, 1.297991173353519e+17, 1.297991173392582e+17, 1.297991173433207e+17, 1.297991173473833e+17, 1.297991173512895e+17, 1.297991173553519e+17, 1.297991173594145e+17, 1.297991173633207e+17, 1.297991173673833e+17, 1.297991173714458e+17, 1.297991173755082e+17, 1.297991173794145e+17, 1.29799117383477e+17, 1.297991173875395e+17, 1.297991173914458e+17, 1.297991173955082e+17, 1.297991173995707e+17, 1.297991174036333e+17, 1.297991174075395e+17, 1.29799117411602e+17, 1.297991174156645e+17, 1.297991174195708e+17, 1.297991174236333e+17, 1.297991174276957e+17, 1.29799117431602e+17, 1.297991174356644e+17, 1.29799117439727e+17, 1.297991174437896e+17, 1.297991174476957e+17, 1.297991174517583e+17, 1.297991174558208e+17, 1.29799117459727e+17, 1.297991174637896e+17, 1.297991174678519e+17, 1.297991174719145e+17, 1.297991174758207e+17, 1.297991174798833e+17, 1.297991174839457e+17, 1.29799117487852e+17, 1.297991174919145e+17, 1.297991174959771e+17, 1.297991174998833e+17, 1.297991175039457e+17, 1.297991175080082e+17, 1.297991175120708e+17, 1.297991175159771e+17, 1.297991175200394e+17, 1.29799117524102e+17, 1.297991175280082e+17, 1.297991175320708e+17, 1.297991175361332e+17, 1.297991175400394e+17, 1.29799117544102e+17, 1.297991175481645e+17, 1.297991175520708e+17, 1.297991175561332e+17, 1.297991175601957e+17, 1.297991175642582e+17, 1.297991175681645e+17, 1.297991175722269e+17, 1.297991175762895e+17, 1.297991175801957e+17, 1.297991175842583e+17, 1.297991175883208e+17, 1.297991175923832e+17, 1.297991175962895e+17, 1.29799117600352e+17, 1.297991176044145e+17, 1.297991176083208e+17, 1.297991176123832e+17, 1.297991176164458e+17, 1.29799117620352e+17, 1.297991176244145e+17, 1.297991176284771e+17, 1.297991176325395e+17, 1.297991176364457e+17, 1.297991176405083e+17, 1.297991176445708e+17, 1.297991176484771e+17, 1.297991176525395e+17, 1.29799117656602e+17, 1.297991176606646e+17, 1.297991176645708e+17, 1.297991176686332e+17, 1.297991176726958e+17, 1.29799117676602e+17, 1.297991176806646e+17, 1.297991176847269e+17, 1.297991176886333e+17, 1.297991176926957e+17, 1.297991176967583e+17, 1.297991177008207e+17, 1.297991177047269e+17, 1.297991177087895e+17, 1.297991177128521e+17, 1.297991177167583e+17, 1.297991177208207e+17, 1.297991177248832e+17, 1.297991177287895e+17, 1.29799117732852e+17, 1.297991177369144e+17, 1.297991177408207e+17, 1.297991177448832e+17, 1.297991177489458e+17, 1.297991177530083e+17, 1.297991177569146e+17, 1.29799117760977e+17, 1.297991177650395e+17, 1.297991177689458e+17, 1.297991177730083e+17, 1.297991177770707e+17, 1.297991177811333e+17, 1.297991177850395e+17, 1.29799117789102e+17, 1.297991177931645e+17, 1.297991177970707e+17, 1.297991178011332e+17, 1.297991178051958e+17, 1.29799117809102e+17, 1.297991178131645e+17, 1.29799117817227e+17, 1.297991178212895e+17, 1.297991178251958e+17, 1.297991178292582e+17, 1.297991178333207e+17, 1.297991178372269e+17, 1.297991178412895e+17, 1.297991178453521e+17, 1.297991178494145e+17, 1.297991178533208e+17, 1.297991178573833e+17, 1.297991178614458e+17, 1.297991178653521e+17, 1.297991178694144e+17, 1.29799117873477e+17, 1.297991178773833e+17, 1.297991178814458e+17, 1.297991178855084e+17, 1.297991178895708e+17, 1.29799117893477e+17, 1.297991178975396e+17, 1.297991179016019e+17, 1.297991179055082e+17, 1.297991179095707e+17, 1.297991179136333e+17, 1.297991179175396e+17, 1.29799117921602e+17, 1.297991179256645e+17, 1.297991179295707e+17, 1.297991179336333e+17, 1.297991179376957e+17, 1.297991179417582e+17, 1.297991179456645e+17, 1.29799117949727e+17, 1.297991179537894e+17, 1.297991179576959e+17, 1.297991179617582e+17, 1.297991179658207e+17, 1.297991179698833e+17, 1.297991179737894e+17, 1.29799117977852e+17, 1.297991179819145e+17, 1.297991179858208e+17, 1.297991179898833e+17, 1.297991179939457e+17, 1.29799117997852e+17, 1.297991180019145e+17, 1.29799118005977e+17, 1.297991180100396e+17, 1.297991180139457e+17, 1.297991180180083e+17, 1.297991180220708e+17, 1.29799118025977e+17, 1.297991180300396e+17, 1.29799118034102e+17, 1.297991180381645e+17, 1.297991180420708e+17, 1.297991180461332e+17, 1.297991180501958e+17, 1.29799118054102e+17, 1.297991180581645e+17, 1.297991180622271e+17, 1.297991180661332e+17, 1.297991180701957e+17, 1.297991180742583e+17, 1.297991180783208e+17, 1.297991180822271e+17, 1.297991180862895e+17, 1.29799118090352e+17, 1.297991180942582e+17, 1.297991180983208e+17, 1.297991181023832e+17, 1.297991181062894e+17, 1.29799118110352e+17, 1.297991181144146e+17, 1.297991181183208e+17, 1.297991181223834e+17, 1.297991181264457e+17, 1.297991181305082e+17, 1.297991181344145e+17, 1.297991181384769e+17, 1.297991181425395e+17, 1.297991181464457e+17, 1.297991181505083e+17, 1.297991181545708e+17, 1.297991181586332e+17, 1.297991181625395e+17, 1.29799118166602e+17, 1.297991181706644e+17, 1.297991181745708e+17, 1.297991181786332e+17, 1.297991181826958e+17, 1.29799118186602e+17, 1.297991181906644e+17, 1.29799118194727e+17, 1.297991181987895e+17, 1.297991182026957e+17, 1.297991182067583e+17, 1.297991182108207e+17, 1.29799118214727e+17, 1.297991182187895e+17, 1.29799118222852e+17, 1.297991182269146e+17, 1.297991182308207e+17, 1.297991182348832e+17, 1.297991182389458e+17, 1.29799118242852e+17, 1.297991182469146e+17, 1.29799118250977e+17, 1.297991182548833e+17, 1.297991182589458e+17, 1.297991182630083e+17, 1.297991182670707e+17, 1.297991182709769e+17, 1.297991182750395e+17, 1.297991182791021e+17, 1.297991182830083e+17, 1.297991182870708e+17, 1.297991182911333e+17, 1.297991182950395e+17, 1.297991182991021e+17, 1.297991183031644e+17, 1.297991183070707e+17, 1.297991183111332e+17, 1.297991183151958e+17, 1.297991183192582e+17, 1.297991183231645e+17, 1.29799118327227e+17, 1.297991183312895e+17, 1.297991183351958e+17, 1.297991183392582e+17, 1.297991183433207e+17, 1.297991183473833e+17, 1.297991183512895e+17, 1.297991183553519e+17, 1.297991183594145e+17, 1.297991183633207e+17, 1.297991183673832e+17, 1.297991183714458e+17, 1.297991183753519e+17, 1.297991183794145e+17, 1.29799118383477e+17, 1.297991183875395e+17, 1.297991183914458e+17, 1.297991183955082e+17, 1.297991183995707e+17, 1.29799118403477e+17, 1.297991184075395e+17, 1.29799118411602e+17, 1.297991184156645e+17, 1.297991184195708e+17, 1.297991184236333e+17, 1.297991184276957e+17, 1.29799118431602e+17, 1.297991184356645e+17, 1.29799118439727e+17, 1.297991184436333e+17, 1.297991184476957e+17, 1.297991184517583e+17, 1.297991184558208e+17, 1.29799118459727e+17, 1.297991184637896e+17, 1.297991184678519e+17, 1.297991184717582e+17, 1.297991184758208e+17, 1.297991184798833e+17, 1.297991184837896e+17, 1.29799118487852e+17, 1.297991184919145e+17, 1.297991184958207e+17, 1.297991184998833e+17, 1.297991185039457e+17, 1.297991185080083e+17, 1.297991185119145e+17, 1.297991185159771e+17, 1.297991185200394e+17, 1.297991185239459e+17, 1.297991185280082e+17, 1.297991185320707e+17, 1.297991185361332e+17, 1.297991185400394e+17, 1.29799118544102e+17, 1.297991185481646e+17, 1.297991185520708e+17, 1.297991185561332e+17, 1.297991185601957e+17, 1.29799118564102e+17, 1.297991185681645e+17, 1.297991185722269e+17, 1.297991185762895e+17, 1.297991185801957e+17, 1.297991185842583e+17, 1.297991185883208e+17, 1.297991185922269e+17, 1.297991185962895e+17, 1.29799118600352e+17, 1.297991186044145e+17, 1.297991186083208e+17, 1.297991186123832e+17, 1.297991186164458e+17, 1.29799118620352e+17, 1.297991186244145e+17, 1.297991186284771e+17, 1.297991186323832e+17, 1.297991186364457e+17, 1.297991186405083e+17, 1.297991186445708e+17, 1.297991186484771e+17, 1.297991186525395e+17, 1.29799118656602e+17, 1.297991186605083e+17, 1.297991186645708e+17},
			             {1.29799100934102e+17, 1.297991009420708e+17, 1.297991009461332e+17, 1.297991009501957e+17, 1.297991009542583e+17, 1.297991009701957e+17},
			             {1.297991015726958e+17, 1.29799101584727e+17, 1.297991015887895e+17},
			             {1.297991016770707e+17, 1.297991016970707e+17},
			             {1.297991017011332e+17, 1.297991017131645e+17},
			             {1.297991017653521e+17, 1.297991017694145e+17, 1.297991017775396e+17, 1.297991017855082e+17, 1.297991017895708e+17},
			             {1.297991017975395e+17, 1.297991018056645e+17},
			             {1.297991018256645e+17, 1.297991018336332e+17},
			             {1.297991018376957e+17, 1.297991018458207e+17},
			             {1.297991019662895e+17, 1.297991019742583e+17},
			             {1.297991019783208e+17, 1.29799101990352e+17},
			             {1.29799102150977e+17, 1.297991021589458e+17},
			             {1.297991021750395e+17, 1.297991021791021e+17},
			             {1.297991022151958e+17, 1.297991022233208e+17},
			             {1.297991022433208e+17, 1.297991022473832e+17},
			             {1.297991024762895e+17, 1.297991024842582e+17},
			             {1.297991024923832e+17, 1.297991025044145e+17, 1.297991025083208e+17, 1.297991025123832e+17},
			             {1.297991025164457e+17, 1.29799102520352e+17, 1.297991025244145e+17, 1.297991025284769e+17},
			             {1.297991025364457e+17, 1.297991025405083e+17, 1.297991025445708e+17, 1.297991025484771e+17},
			             {1.297991025967583e+17, 1.297991026008207e+17, 1.297991026087895e+17},
			             {1.297991026931644e+17, 1.297991027131645e+17},
			             {1.297991028095708e+17, 1.297991028256645e+17, 1.297991028295708e+17, 1.297991028376957e+17, 1.297991028456645e+17},
			             {1.29799102905977e+17, 1.297991029220708e+17},
			             {1.297991029381645e+17, 1.297991029461332e+17, 1.297991029501957e+17},
			             {1.29799117242852e+17, 1.297991172951958e+17},
			             {1.297991060664458e+17, 1.297991060705083e+17, 1.297991060786333e+17, 1.29799106086602e+17, 1.297991060945708e+17},
			             {1.297991062953521e+17, 1.29799106303477e+17, 1.297991063075396e+17, 1.297991063155084e+17, 1.297991063195707e+17, 1.29799106323477e+17, 1.297991063275396e+17, 1.297991063316019e+17, 1.297991063356645e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}}, {{}, {}, {}}, {{}, {}}, {{}, {}}, {{}, {}, {}, {}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}, {}, {}}, {{}, {}, {}, {}}, {{}, {}, {}, {}}, {{}, {}, {}}, {{}, {}}, {{}, {}, {}, {}, {}}, {{}, {}}, {{}, {}, {}}, {{}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
