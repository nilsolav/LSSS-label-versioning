netcdf mask {
	:date_created = "20200810T140900";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200810T140900";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 1;
			channels = 6;
			categories = 6;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0;
			max_depth =  53.5;
			start_time = 131381777062669440;
			end_time = 131381784329544448;
			region_id = 1;
			region_name = "Layer1";
			region_provenance = "LSSS";
			region_comment = "";
			region_category_names = "0", "0", "0", "0", "0", "0";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1, 2, 3, 4, 5, 6;
			region_type = analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63;
			mask_times = {1.313817770626694e+17, 1.313817770695446e+17, 1.313817770718883e+17, 1.313817770832945e+17, 1.313817770865757e+17, 1.313817770934508e+17, 1.313817770997007e+17, 1.313817771045445e+17, 1.313817771139195e+17, 1.31381777117982e+17, 1.313817771239195e+17, 1.313817771314195e+17, 1.313817771384508e+17, 1.313817771450132e+17, 1.313817771534508e+17, 1.313817771582945e+17, 1.313817771662633e+17, 1.313817771751695e+17, 1.313817771797007e+17, 1.31381777186107e+17, 1.313817771925133e+17, 1.313817771995444e+17, 1.313817772062633e+17, 1.31381777208607e+17, 1.313817772201696e+17, 1.313817772225133e+17, 1.31381777224857e+17, 1.313817772365757e+17, 1.313817772389196e+17, 1.31381777246732e+17, 1.313817772528257e+17, 1.313817772595444e+17, 1.31381777266107e+17, 1.31381777272982e+17, 1.313817772797007e+17, 1.313817772865757e+17, 1.313817772931383e+17, 1.313817773001695e+17, 1.313817773065757e+17, 1.313817773137633e+17, 1.31381777319857e+17, 1.31381777326732e+17, 1.313817773337633e+17, 1.313817773406382e+17, 1.313817773473569e+17, 1.313817773542319e+17, 1.31381777360482e+17, 1.313817773678258e+17, 1.313817773742319e+17, 1.313817773811071e+17, 1.313817773895444e+17, 1.313817773931382e+17, 1.313817773993883e+17, 1.313817774057944e+17, 1.313817774118883e+17, 1.31381777418607e+17, 1.313817774256383e+17, 1.313817774312632e+17, 1.313817774375132e+17, 1.313817774445445e+17, 1.313817774468883e+17, 1.313817774587633e+17, 1.313817774628257e+17, 1.313817774651695e+17, 1.313817774770445e+17, 1.313817774814195e+17, 1.313817774837633e+17, 1.313817774950132e+17, 1.313817774993883e+17, 1.31381777506107e+17, 1.31381777513607e+17, 1.313817775187633e+17, 1.313817775276695e+17, 1.313817775326696e+17, 1.313817775422008e+17, 1.313817775457946e+17, 1.313817775526694e+17, 1.313817775584507e+17, 1.313817775645445e+17, 1.31381777571732e+17, 1.313817775784507e+17, 1.313817775853257e+17, 1.313817775918883e+17, 1.313817775981382e+17, 1.313817776042321e+17, 1.313817776111069e+17, 1.313817776181382e+17, 1.313817776251695e+17, 1.313817776311069e+17, 1.313817776375133e+17, 1.313817776454821e+17, 1.313817776511071e+17, 1.313817776565757e+17, 1.313817776640756e+17, 1.313817776707945e+17, 1.313817776768882e+17, 1.313817776851695e+17, 1.313817776887633e+17, 1.313817776962632e+17, 1.31381777701732e+17, 1.313817777100132e+17, 1.313817777168882e+17, 1.313817777211069e+17, 1.313817777281382e+17, 1.313817777350132e+17, 1.313817777412632e+17, 1.31381777747982e+17, 1.31381777752357e+17, 1.313817777611071e+17, 1.313817777678258e+17, 1.313817777745445e+17, 1.313817777806382e+17, 1.313817777875132e+17, 1.313817777943884e+17, 1.313817778062632e+17, 1.313817778098569e+17, 1.313817778168883e+17, 1.313817778228257e+17, 1.313817778295444e+17, 1.31381777836107e+17, 1.313817778425133e+17, 1.313817778495446e+17, 1.313817778518883e+17, 1.313817778600133e+17, 1.313817778645444e+17, 1.313817778726696e+17, 1.313817778772008e+17, 1.313817778840758e+17, 1.313817778909508e+17, 1.313817778972008e+17, 1.313817779040756e+17, 1.313817779101695e+17, 1.313817779170445e+17, 1.31381777923607e+17, 1.31381777930482e+17, 1.313817779328257e+17, 1.313817779443884e+17, 1.313817779482945e+17, 1.313817779568882e+17, 1.31381777959232e+17, 1.313817779684507e+17, 1.313817779725133e+17, 1.313817779784508e+17, 1.313817779851695e+17, 1.313817779937632e+17, 1.313817779972008e+17, 1.313817780057946e+17, 1.31381778009857e+17, 1.31381778016732e+17, 1.313817780236069e+17, 1.313817780306383e+17, 1.313817780426696e+17, 1.313817780453257e+17, 1.313817780507945e+17, 1.313817780579821e+17, 1.313817780632945e+17, 1.313817780700133e+17, 1.31381778072357e+17, 1.313817780843882e+17, 1.31381778086732e+17, 1.313817780984507e+17, 1.313817781007945e+17, 1.31381778108607e+17, 1.313817781181382e+17, 1.31381778120482e+17, 1.313817781276695e+17, 1.313817781339196e+17, 1.313817781417321e+17, 1.313817781487633e+17, 1.31381778155482e+17, 1.313817781626696e+17, 1.313817781725132e+17, 1.31381778174857e+17, 1.313817781814195e+17, 1.313817781859507e+17, 1.313817781925133e+17, 1.313817781993883e+17, 1.313817782059507e+17, 1.313817782082945e+17, 1.31381778219857e+17, 1.313817782251695e+17, 1.313817782318883e+17, 1.313817782387633e+17, 1.313817782411069e+17, 1.313817782525133e+17, 1.313817782568882e+17, 1.313817782603258e+17, 1.31381778270482e+17, 1.313817782770445e+17, 1.313817782859507e+17, 1.313817782911069e+17, 1.313817782932945e+17, 1.313817783018883e+17, 1.313817783115757e+17, 1.313817783156383e+17, 1.313817783179821e+17, 1.313817783295446e+17, 1.313817783318883e+17, 1.313817783428257e+17, 1.31381778345482e+17, 1.313817783532945e+17, 1.31381778356107e+17, 1.313817783637632e+17, 1.313817783673571e+17, 1.313817783747008e+17, 1.313817783815757e+17, 1.313817783884508e+17, 1.313817783953257e+17, 1.313817784018883e+17, 1.313817784081382e+17, 1.313817784150132e+17, 1.313817784257944e+17, 1.313817784290757e+17, 1.313817784345445e+17, 1.313817784422007e+17, 1.313817784470445e+17, 1.313817784542321e+17, 1.313817784628257e+17, 1.313817784679821e+17, 1.313817784797007e+17, 1.313817784820445e+17, 1.313817784857946e+17, 1.313817784945444e+17, 1.313817785042319e+17, 1.313817785065757e+17, 1.31381778512982e+17, 1.313817785178258e+17, 1.313817785273569e+17, 1.313817785326696e+17, 1.313817785415758e+17, 1.313817785443882e+17, 1.31381778551732e+17, 1.313817785540756e+17, 1.313817785640758e+17, 1.313817785664196e+17, 1.31381778576107e+17, 1.313817785784507e+17, 1.313817785889196e+17, 1.313817785939195e+17, 1.313817786011071e+17, 1.313817786081382e+17, 1.313817786151695e+17, 1.313817786207945e+17, 1.313817786278258e+17, 1.313817786301696e+17, 1.313817786372008e+17, 1.313817786434508e+17, 1.31381778649232e+17, 1.31381778655482e+17, 1.313817786639195e+17, 1.313817786675132e+17, 1.31381778675482e+17, 1.31381778679232e+17, 1.313817786859507e+17, 1.313817786925132e+17, 1.313817786982945e+17, 1.313817787050132e+17, 1.313817787109508e+17, 1.313817787181382e+17, 1.31381778724857e+17, 1.313817787315758e+17, 1.313817787384508e+17, 1.313817787451695e+17, 1.313817787520444e+17, 1.313817787581382e+17, 1.313817787656383e+17, 1.313817787725133e+17, 1.313817787806382e+17, 1.313817787873569e+17, 1.313817787931383e+17, 1.313817788000133e+17, 1.313817788114195e+17, 1.313817788137632e+17, 1.313817788193883e+17, 1.313817788245445e+17, 1.313817788270445e+17, 1.313817788384507e+17, 1.313817788412632e+17, 1.313817788504819e+17, 1.313817788543882e+17, 1.31381778860482e+17, 1.313817788662632e+17, 1.313817788739195e+17, 1.313817788807945e+17, 1.313817788876695e+17, 1.313817788939195e+17, 1.313817789006382e+17, 1.313817789072008e+17, 1.313817789143882e+17, 1.313817789206383e+17, 1.313817789275132e+17, 1.31381778933607e+17, 1.313817789403258e+17, 1.313817789464195e+17, 1.313817789534508e+17, 1.313817789603258e+17, 1.313817789672006e+17, 1.313817789731383e+17, 1.31381778979857e+17, 1.313817789822007e+17, 1.313817789889196e+17, 1.313817789942321e+17, 1.313817790039195e+17, 1.313817790097007e+17, 1.313817790165757e+17, 1.313817790189196e+17, 1.313817790303256e+17, 1.313817790342321e+17, 1.313817790415757e+17, 1.313817790472008e+17, 1.313817790547007e+17, 1.313817790601695e+17, 1.313817790675132e+17, 1.313817790750132e+17, 1.313817790801695e+17, 1.313817790868882e+17, 1.313817790932945e+17, 1.313817790995444e+17, 1.313817791070445e+17, 1.313817791137633e+17, 1.313817791207945e+17, 1.31381779130482e+17, 1.313817791347007e+17, 1.313817791406383e+17, 1.313817791465757e+17, 1.313817791532945e+17, 1.313817791589196e+17, 1.313817791695444e+17, 1.313817791718883e+17, 1.31381779179857e+17, 1.313817791853257e+17, 1.313817791932945e+17, 1.313817792022007e+17, 1.31381779206107e+17, 1.313817792120444e+17, 1.313817792184508e+17, 1.31381779224857e+17, 1.313817792314195e+17, 1.31381779237982e+17, 1.313817792447007e+17, 1.313817792511071e+17, 1.313817792576695e+17, 1.31381779264857e+17, 1.313817792703258e+17, 1.313817792770445e+17, 1.313817792842319e+17, 1.313817792925133e+17, 1.313817792972008e+17, 1.313817793031382e+17, 1.313817793101695e+17, 1.313817793187633e+17, 1.313817793232945e+17, 1.313817793307945e+17, 1.31381779335482e+17, 1.313817793415758e+17, 1.313817793501695e+17, 1.313817793547007e+17, 1.313817793628259e+17, 1.313817793689196e+17, 1.313817793773571e+17, 1.313817793820444e+17, 1.313817793843882e+17, 1.31381779396107e+17, 1.313817794020444e+17, 1.313817794078258e+17, 1.31381779419232e+17, 1.313817794217321e+17, 1.31381779428607e+17, 1.31381779435482e+17, 1.313817794425133e+17, 1.31381779449232e+17, 1.313817794545445e+17, 1.313817794625133e+17, 1.31381779468607e+17, 1.313817794773571e+17, 1.313817794806383e+17, 1.313817794882944e+17, 1.313817794943882e+17, 1.313817795034508e+17, 1.313817795095444e+17, 1.313817795170445e+17, 1.313817795250132e+17, 1.313817795365757e+17, 1.31381779539232e+17, 1.313817795500133e+17, 1.313817795528257e+17, 1.313817795601695e+17, 1.313817795662633e+17, 1.313817795742321e+17, 1.313817795812632e+17, 1.313817795881382e+17, 1.313817795959507e+17, 1.313817796031383e+17, 1.313817796107945e+17, 1.31381779618607e+17, 1.31381779625482e+17, 1.31381779632357e+17, 1.313817796347008e+17, 1.31381779646732e+17, 1.313817796507945e+17, 1.313817796607945e+17, 1.31381779664857e+17, 1.313817796753257e+17, 1.313817796778257e+17, 1.313817796887633e+17, 1.313817796911071e+17, 1.313817796978258e+17, 1.313817797001695e+17, 1.313817797106382e+17, 1.313817797142321e+17, 1.313817797220445e+17, 1.313817797243884e+17, 1.313817797359507e+17, 1.31381779738607e+17, 1.313817797492321e+17, 1.313817797520444e+17, 1.31381779757982e+17, 1.313817797653257e+17, 1.313817797734508e+17, 1.313817797803258e+17, 1.313817797870445e+17, 1.313817797939195e+17, 1.313817798009508e+17, 1.313817798073569e+17, 1.313817798137632e+17, 1.313817798206382e+17, 1.313817798270445e+17, 1.313817798293883e+17, 1.313817798407945e+17, 1.313817798451695e+17, 1.313817798522007e+17, 1.313817798590757e+17, 1.313817798657946e+17, 1.313817798731383e+17, 1.313817798784507e+17, 1.313817798853257e+17, 1.31381779892357e+17, 1.313817798947008e+17, 1.313817799062632e+17, 1.313817799134508e+17, 1.313817799187633e+17, 1.313817799259508e+17, 1.313817799351695e+17, 1.31381779939232e+17, 1.313817799481382e+17, 1.313817799531382e+17, 1.313817799603258e+17, 1.313817799668883e+17, 1.313817799732945e+17, 1.313817799804819e+17, 1.313817799882945e+17, 1.313817799925133e+17, 1.313817799981382e+17, 1.313817800064195e+17, 1.313817800137632e+17, 1.313817800193883e+17, 1.31381780021732e+17, 1.313817800240756e+17, 1.31381780026732e+17, 1.31381780029857e+17, 1.313817800323571e+17, 1.313817800456383e+17, 1.313817800493883e+17, 1.313817800557944e+17, 1.313817800620445e+17, 1.31381780068607e+17, 1.313817800762633e+17, 1.313817800809508e+17, 1.313817800872008e+17, 1.313817800940756e+17, 1.313817801018883e+17, 1.313817801095446e+17, 1.313817801170445e+17, 1.313817801237632e+17, 1.313817801312632e+17, 1.313817801382945e+17, 1.31381780144857e+17, 1.313817801522007e+17, 1.31381780159857e+17, 1.313817801622007e+17, 1.313817801693883e+17, 1.31381780171732e+17, 1.313817801750132e+17, 1.313817801775133e+17, 1.313817801801695e+17, 1.313817801825133e+17, 1.313817801875132e+17, 1.313817801900132e+17, 1.313817801934508e+17, 1.313817801973569e+17, 1.31381780199857e+17, 1.31381780209857e+17, 1.31381780212357e+17, 1.313817802187633e+17, 1.313817802212634e+17, 1.31381780226107e+17, 1.313817802315758e+17, 1.313817802340758e+17, 1.31381780237982e+17, 1.313817802439195e+17, 1.313817802476695e+17, 1.31381780254857e+17, 1.313817802593882e+17, 1.313817802664196e+17, 1.313817802722007e+17, 1.31381780277982e+17, 1.313817802837633e+17, 1.313817802903256e+17, 1.313817802959508e+17, 1.313817803028257e+17, 1.313817803078257e+17, 1.313817803131383e+17, 1.31381780317982e+17, 1.31381780322357e+17, 1.313817803275133e+17, 1.313817803326694e+17, 1.313817803378258e+17, 1.313817803447008e+17, 1.313817803504819e+17, 1.313817803528257e+17, 1.313817803551695e+17, 1.313817803576695e+17, 1.313817803609508e+17, 1.313817803642319e+17, 1.31381780366732e+17, 1.313817803770445e+17, 1.31381780379857e+17, 1.313817803822008e+17, 1.31381780389232e+17, 1.313817803926696e+17, 1.313817803987633e+17, 1.313817804031382e+17, 1.313817804081382e+17, 1.313817804128257e+17, 1.31381780418607e+17, 1.313817804228257e+17, 1.31381780427982e+17, 1.313817804334508e+17, 1.313817804357944e+17, 1.313817804428257e+17, 1.31381780448607e+17, 1.313817804534508e+17, 1.31381780459232e+17, 1.313817804628257e+17, 1.313817804681382e+17, 1.313817804731382e+17, 1.31381780478607e+17, 1.313817804828257e+17, 1.313817804886071e+17, 1.313817804925133e+17, 1.313817805065757e+17, 1.313817805122008e+17, 1.313817805197007e+17, 1.313817805265757e+17, 1.31381780532357e+17, 1.313817805395446e+17, 1.313817805473569e+17, 1.313817805532945e+17, 1.313817805590758e+17, 1.313817805659507e+17, 1.31381780570482e+17, 1.31381780579857e+17, 1.313817805822008e+17, 1.313817805940756e+17, 1.313817805964195e+17, 1.31381780607982e+17, 1.313817806103258e+17, 1.31381780618607e+17, 1.313817806231382e+17, 1.313817806309508e+17, 1.313817806389194e+17, 1.313817806456383e+17, 1.313817806543884e+17, 1.313817806568883e+17, 1.313817806670445e+17, 1.313817806726696e+17, 1.313817806815757e+17, 1.313817806872008e+17, 1.313817806951695e+17, 1.313817807020444e+17, 1.313817807090758e+17, 1.313817807170445e+17, 1.313817807225133e+17, 1.31381780729232e+17, 1.313817807315758e+17, 1.31381780743607e+17, 1.313817807459507e+17, 1.31381780755482e+17, 1.31381780759857e+17, 1.313817807622007e+17, 1.31381780774857e+17, 1.313817807807945e+17, 1.313817807872008e+17, 1.313817807942321e+17, 1.313817808001696e+17, 1.313817808068883e+17, 1.31381780809232e+17, 1.313817808206382e+17, 1.313817808231382e+17, 1.313817808328257e+17, 1.313817808351694e+17, 1.313817808462633e+17, 1.31381780851732e+17, 1.313817808590758e+17, 1.313817808614195e+17, 1.313817808732945e+17, 1.313817808756383e+17, 1.31381780884857e+17, 1.313817808890757e+17, 1.313817808959507e+17, 1.31381780902982e+17, 1.313817809101695e+17, 1.31381780916732e+17, 1.313817809239195e+17, 1.313817809306382e+17, 1.313817809375133e+17, 1.313817809434508e+17, 1.31381780950482e+17, 1.31381780959232e+17, 1.313817809634508e+17, 1.313817809700132e+17, 1.313817809767319e+17, 1.313817809848571e+17, 1.313817809872008e+17, 1.313817810009508e+17, 1.313817810032945e+17, 1.313817810111071e+17, 1.313817810134508e+17, 1.313817810253257e+17, 1.313817810276695e+17, 1.313817810339195e+17, 1.313817810412632e+17, 1.313817810482944e+17, 1.31381781059857e+17, 1.313817810632946e+17, 1.313817810717321e+17, 1.31381781076107e+17, 1.313817810832945e+17, 1.313817810889196e+17, 1.313817810956383e+17, 1.313817810984508e+17, 1.31381781103607e+17, 1.313817811101696e+17, 1.313817811170445e+17, 1.313817811242321e+17, 1.31381781132357e+17, 1.313817811431382e+17, 1.313817811462633e+17, 1.313817811542319e+17, 1.313817811586071e+17, 1.313817811668882e+17, 1.313817811757944e+17, 1.313817811809507e+17, 1.313817811879821e+17, 1.313817811940758e+17, 1.313817812012632e+17, 1.313817812128257e+17, 1.313817812151695e+17, 1.31381781222357e+17, 1.313817812268883e+17, 1.313817812331382e+17, 1.31381781239857e+17, 1.313817812497007e+17, 1.313817812550132e+17, 1.313817812626694e+17, 1.313817812697007e+17, 1.313817812728257e+17, 1.313817812845445e+17, 1.313817812909508e+17, 1.313817813011069e+17, 1.313817813064196e+17, 1.31381781312982e+17, 1.313817813153258e+17, 1.31381781326732e+17, 1.313817813290757e+17, 1.313817813372008e+17, 1.313817813420445e+17, 1.313817813500133e+17, 1.313817813573571e+17, 1.313817813672008e+17, 1.313817813707945e+17, 1.313817813776695e+17, 1.313817813839195e+17, 1.313817813862632e+17, 1.313817813979821e+17, 1.313817814022008e+17, 1.313817814122007e+17, 1.313817814145445e+17, 1.313817814209508e+17, 1.313817814257944e+17, 1.313817814315758e+17, 1.313817814373569e+17, 1.31381781446107e+17, 1.313817814509508e+17, 1.313817814573569e+17, 1.31381781463607e+17, 1.313817814700132e+17, 1.313817814757946e+17, 1.313817814834508e+17, 1.313817814893883e+17, 1.313817814965757e+17, 1.313817815056383e+17, 1.313817815090757e+17, 1.31381781516732e+17, 1.313817815215757e+17, 1.313817815275133e+17, 1.313817815347008e+17, 1.313817815436069e+17, 1.313817815487633e+17, 1.313817815551695e+17, 1.313817815618883e+17, 1.313817815695444e+17, 1.313817815747008e+17, 1.313817815803258e+17, 1.313817815872008e+17, 1.313817815943882e+17, 1.313817816012632e+17, 1.313817816073569e+17, 1.313817816145445e+17, 1.313817816207945e+17, 1.313817816276695e+17, 1.313817816348571e+17, 1.313817816415758e+17, 1.313817816478258e+17, 1.31381781655482e+17, 1.31381781663607e+17, 1.313817816687631e+17, 1.31381781676732e+17, 1.313817816839195e+17, 1.313817816918883e+17, 1.313817816978257e+17, 1.31381781705482e+17, 1.313817817134508e+17, 1.313817817206383e+17, 1.313817817275132e+17, 1.313817817350132e+17, 1.313817817418883e+17, 1.313817817482944e+17, 1.31381781755482e+17, 1.313817817614195e+17, 1.313817817714194e+17, 1.313817817739195e+17, 1.313817817804819e+17, 1.313817817828257e+17, 1.313817817931383e+17, 1.313817817972008e+17, 1.31381781804857e+17, 1.313817818103258e+17, 1.313817818175132e+17, 1.31381781822982e+17, 1.31381781829857e+17, 1.313817818378258e+17, 1.313817818443882e+17, 1.313817818495444e+17, 1.313817818581382e+17, 1.313817818667319e+17, 1.313817818714195e+17, 1.313817818773571e+17, 1.313817818845445e+17, 1.313817818907945e+17, 1.313817818978257e+17, 1.313817819047008e+17, 1.313817819115757e+17, 1.313817819175132e+17, 1.313817819247008e+17, 1.313817819318883e+17, 1.313817819390757e+17, 1.313817819456383e+17, 1.313817819525133e+17, 1.313817819643882e+17, 1.31381781966732e+17, 1.313817819747008e+17, 1.31381781982982e+17, 1.313817819926696e+17, 1.313817819950132e+17, 1.31381782002357e+17, 1.313817820084508e+17, 1.31381782014857e+17, 1.31381782021732e+17, 1.313817820339195e+17, 1.313817820362633e+17, 1.313817820432945e+17, 1.313817820489194e+17, 1.313817820597007e+17, 1.313817820622008e+17, 1.313817820687633e+17, 1.313817820751695e+17, 1.313817820828257e+17, 1.313817820890757e+17, 1.313817820959507e+17, 1.313817821020445e+17, 1.31381782109232e+17, 1.313817821157944e+17, 1.31381782122982e+17, 1.31381782129857e+17, 1.313817821387633e+17, 1.313817821451695e+17, 1.313817821514195e+17, 1.313817821586071e+17, 1.31381782165482e+17, 1.313817821725133e+17, 1.313817821787633e+17, 1.313817821856383e+17, 1.31381782192357e+17, 1.313817821993883e+17, 1.313817822059508e+17, 1.313817822131382e+17, 1.31381782216107e+17, 1.313817822268883e+17, 1.313817822357946e+17, 1.313817822381382e+17, 1.313817822406383e+17, 1.31381782242982e+17, 1.313817822557946e+17, 1.313817822614195e+17, 1.313817822682944e+17, 1.313817822751695e+17, 1.313817822811069e+17, 1.313817822918883e+17, 1.313817822953257e+17, 1.313817823020445e+17, 1.313817823084507e+17, 1.313817823259507e+17, 1.313817823300133e+17, 1.31381782339232e+17, 1.313817823462633e+17, 1.313817823534508e+17, 1.313817823593883e+17, 1.313817823673569e+17, 1.31381782372982e+17, 1.313817823800132e+17, 1.313817823868882e+17, 1.313817823937633e+17, 1.313817823993883e+17, 1.313817824059507e+17, 1.313817824082945e+17, 1.313817824200132e+17, 1.313817824243882e+17, 1.313817824329819e+17, 1.313817824400133e+17, 1.313817824468882e+17, 1.313817824531383e+17, 1.31381782460482e+17, 1.313817824670445e+17, 1.313817824742319e+17, 1.313817824765757e+17, 1.313817824889194e+17, 1.313817824950132e+17, 1.313817825022007e+17, 1.313817825093883e+17, 1.313817825156383e+17, 1.313817825226694e+17, 1.313817825293883e+17, 1.313817825364196e+17, 1.313817825418883e+17, 1.313817825487633e+17, 1.313817825557946e+17, 1.313817825628257e+17, 1.313817825725133e+17, 1.31381782576107e+17, 1.313817825822008e+17, 1.313817825890757e+17, 1.313817825959508e+17, 1.31381782602982e+17, 1.313817826095444e+17, 1.313817826162633e+17, 1.313817826231382e+17, 1.313817826300133e+17, 1.31381782636732e+17, 1.313817826440758e+17, 1.313817826509508e+17, 1.313817826575132e+17, 1.313817826645445e+17, 1.31381782671732e+17, 1.313817826797007e+17, 1.313817826887633e+17, 1.313817826940756e+17, 1.313817826964195e+17, 1.313817827095446e+17, 1.313817827128257e+17, 1.313817827197007e+17, 1.313817827259508e+17, 1.31381782731732e+17, 1.313817827387633e+17, 1.313817827459507e+17, 1.313817827531382e+17, 1.313817827606383e+17, 1.313817827675132e+17, 1.313817827753257e+17, 1.313817827826694e+17, 1.313817827906382e+17, 1.313817827951695e+17, 1.31381782802357e+17, 1.313817828047007e+17, 1.313817828164195e+17, 1.313817828220445e+17, 1.313817828301695e+17, 1.313817828372008e+17, 1.313817828439196e+17, 1.313817828500133e+17, 1.313817828570445e+17, 1.313817828650132e+17, 1.313817828675133e+17, 1.313817828815758e+17, 1.313817828840758e+17, 1.313817828926694e+17, 1.313817828970445e+17, 1.31381782903607e+17, 1.313817829134508e+17, 1.31381782920482e+17, 1.313817829332945e+17, 1.313817829356383e+17, 1.313817829379821e+17, 1.313817829411071e+17, 1.313817829434508e+17, 1.313817829457944e+17, 1.313817829481382e+17, 1.31381782951732e+17, 1.313817829539195e+17, 1.313817829562633e+17, 1.313817829584507e+17, 1.313817829607945e+17, 1.31381782962982e+17, 1.313817829651695e+17, 1.313817829675132e+17, 1.313817829697007e+17, 1.313817829720445e+17, 1.313817829743882e+17, 1.313817829765757e+17, 1.313817829789196e+17, 1.313817829811071e+17, 1.313817829834508e+17, 1.313817829856383e+17, 1.31381782987982e+17, 1.313817829901695e+17, 1.31381782992357e+17, 1.313817829956383e+17, 1.313817829978258e+17, 1.313817830003256e+17, 1.313817830025133e+17, 1.313817830047007e+17, 1.313817830070445e+17, 1.313817830101695e+17, 1.31381783012357e+17, 1.313817830145445e+17, 1.313817830176695e+17, 1.313817830200133e+17, 1.313817830222007e+17, 1.313817830245445e+17, 1.31381783026732e+17, 1.313817830290757e+17, 1.313817830314195e+17, 1.31381783033607e+17, 1.313817830359507e+17, 1.313817830382945e+17, 1.313817830404819e+17, 1.313817830428257e+17, 1.313817830450132e+17, 1.313817830472006e+17, 1.313817830503258e+17, 1.313817830526694e+17, 1.313817830550132e+17, 1.313817830572008e+17, 1.313817830595444e+17, 1.31381783061732e+17, 1.313817830640756e+17, 1.313817830662633e+17, 1.313817830686071e+17, 1.313817830707945e+17, 1.31381783072982e+17, 1.313817830753257e+17, 1.313817830775132e+17, 1.31381783079857e+17, 1.31381783082982e+17, 1.313817830853257e+17, 1.313817830875133e+17, 1.31381783089857e+17, 1.313817830920444e+17, 1.313817830943882e+17, 1.313817830965757e+17, 1.313817830987633e+17, 1.313817831011071e+17, 1.313817831032946e+17, 1.313817831056383e+17, 1.313817831078257e+17, 1.313817831101695e+17, 1.313817831123571e+17, 1.313817831145445e+17, 1.313817831168883e+17, 1.31381783119232e+17, 1.313817831215757e+17, 1.313817831237632e+17, 1.313817831267319e+17, 1.313817831290757e+17, 1.313817831314195e+17, 1.31381783133607e+17, 1.313817831359507e+17, 1.313817831381382e+17, 1.313817831403258e+17, 1.313817831426696e+17, 1.31381783144857e+17, 1.313817831472008e+17, 1.313817831493883e+17, 1.31381783151732e+17, 1.313817831539195e+17, 1.313817831562633e+17, 1.313817831593883e+17, 1.31381783161732e+17, 1.313817831639195e+17, 1.31381783166107e+17, 1.313817831684507e+17, 1.313817831706383e+17, 1.31381783172982e+17, 1.313817831751695e+17, 1.313817831775132e+17, 1.313817831797007e+17, 1.313817831820444e+17, 1.313817831842319e+17, 1.313817831864196e+17, 1.313817831887633e+17, 1.313817831909508e+17, 1.313817831932945e+17, 1.313817831956383e+17, 1.313817831978257e+17, 1.313817832001695e+17, 1.313817832032945e+17, 1.313817832056383e+17, 1.313817832078258e+17, 1.313817832101696e+17, 1.31381783212357e+17, 1.313817832147007e+17, 1.313817832168883e+17, 1.31381783219232e+17, 1.313817832215757e+17, 1.313817832237632e+17, 1.313817832259508e+17, 1.313817832282945e+17, 1.313817832304819e+17, 1.313817832328257e+17, 1.313817832359507e+17, 1.313817832382945e+17, 1.313817832406382e+17, 1.313817832428257e+17, 1.313817832451694e+17, 1.313817832473571e+17, 1.313817832497007e+17, 1.313817832518883e+17, 1.313817832542319e+17, 1.313817832564196e+17, 1.31381783258607e+17, 1.313817832609507e+17, 1.313817832631383e+17, 1.31381783265482e+17, 1.313817832686071e+17, 1.313817832709508e+17, 1.313817832731382e+17, 1.31381783275482e+17, 1.313817832778257e+17, 1.313817832800133e+17, 1.31381783282357e+17, 1.313817832845445e+17, 1.313817832875132e+17, 1.313817832906382e+17, 1.313817832928257e+17, 1.313817832950132e+17, 1.313817832973571e+17, 1.313817832995446e+17, 1.313817833018883e+17, 1.313817833040758e+17, 1.313817833064195e+17, 1.313817833086071e+17, 1.313817833109508e+17, 1.313817833131383e+17, 1.313817833153258e+17, 1.313817833176695e+17, 1.31381783319857e+17, 1.313817833222007e+17, 1.313817833243884e+17, 1.31381783326732e+17, 1.313817833289196e+17, 1.313817833311071e+17, 1.313817833342321e+17, 1.313817833365757e+17, 1.313817833387633e+17, 1.313817833411069e+17, 1.313817833432945e+17, 1.313817833456383e+17, 1.313817833478257e+17, 1.313817833501695e+17, 1.31381783352357e+17, 1.313817833545444e+17, 1.313817833568882e+17, 1.31381783359232e+17, 1.313817833614195e+17, 1.313817833637632e+17, 1.313817833668883e+17, 1.313817833693883e+17, 1.313817833715757e+17, 1.313817833737632e+17, 1.31381783376107e+17, 1.313817833782944e+17, 1.313817833806382e+17, 1.313817833828257e+17, 1.313817833851695e+17, 1.313817833875132e+17, 1.313817833897007e+17, 1.313817833920445e+17, 1.313817833942321e+17, 1.313817833965757e+17, 1.313817833997007e+17, 1.313817834020445e+17, 1.313817834042319e+17, 1.313817834064196e+17, 1.313817834087633e+17, 1.313817834109508e+17, 1.313817834132945e+17, 1.313817834156383e+17, 1.313817834178258e+17, 1.313817834201695e+17, 1.31381783422357e+17, 1.313817834247008e+17, 1.313817834270446e+17, 1.31381783429232e+17, 1.313817834325133e+17, 1.313817834347007e+17, 1.313817834370445e+17, 1.31381783439232e+17, 1.313817834415758e+17, 1.313817834437632e+17, 1.313817834459507e+17, 1.313817834482945e+17, 1.313817834504819e+17, 1.313817834528257e+17, 1.313817834550132e+17, 1.313817834573571e+17, 1.313817834595444e+17, 1.31381783461732e+17, 1.313817834640758e+17, 1.313817834662632e+17, 1.31381783468607e+17, 1.313817834707945e+17, 1.313817834731383e+17, 1.313817834762633e+17, 1.313817834784507e+17, 1.313817834806383e+17, 1.31381783482982e+17, 1.313817834851695e+17, 1.313817834875132e+17, 1.313817834897009e+17, 1.313817834920445e+17, 1.313817834942319e+17, 1.313817834965757e+17, 1.313817834987633e+17, 1.313817835009508e+17, 1.313817835032945e+17, 1.313817835054821e+17, 1.31381783508607e+17, 1.313817835109508e+17, 1.313817835132946e+17, 1.313817835156383e+17, 1.313817835178258e+17, 1.313817835201695e+17, 1.31381783522357e+17, 1.313817835256383e+17, 1.313817835279821e+17, 1.313817835307945e+17, 1.313817835331382e+17, 1.313817835362632e+17, 1.31381783538607e+17, 1.31381783541732e+17, 1.313817835439195e+17, 1.313817835462633e+17, 1.313817835484507e+17, 1.313817835507944e+17, 1.31381783552982e+17, 1.313817835551695e+17, 1.313817835575132e+17, 1.313817835597007e+17, 1.313817835620445e+17, 1.313817835642319e+17, 1.313817835665756e+17, 1.313817835687633e+17, 1.313817835709508e+17, 1.313817835737632e+17, 1.313817835759508e+17, 1.313817835782945e+17, 1.31381783580482e+17, 1.313817835828257e+17, 1.313817835853257e+17, 1.313817835876695e+17, 1.31381783589857e+17, 1.313817835922007e+17, 1.313817835943882e+17, 1.31381783596732e+17, 1.313817835989196e+17, 1.313817836012632e+17, 1.313817836034508e+17, 1.313817836057946e+17, 1.31381783607982e+17, 1.313817836101695e+17, 1.313817836125133e+17, 1.313817836147008e+17, 1.31381783617982e+17, 1.313817836201695e+17, 1.313817836225132e+17, 1.31381783624857e+17, 1.313817836270445e+17, 1.313817836293883e+17, 1.313817836315757e+17, 1.313817836339195e+17, 1.31381783636107e+17, 1.313817836384508e+17, 1.313817836406382e+17, 1.313817836428257e+17, 1.313817836451695e+17, 1.313817836473569e+17, 1.313817836497007e+17, 1.313817836518883e+17, 1.313817836542321e+17, 1.313817836564195e+17, 1.313817836587633e+17, 1.31381783661732e+17, 1.313817836640758e+17, 1.313817836662632e+17, 1.31381783668607e+17, 1.313817836707945e+17, 1.313817836731383e+17, 1.313817836753257e+17, 1.313817836776695e+17, 1.313817836800132e+17, 1.313817836822008e+17, 1.313817836845445e+17, 1.31381783686732e+17, 1.313817836890757e+17, 1.313817836912632e+17, 1.313817836943884e+17, 1.31381783696732e+17, 1.313817836989196e+17, 1.313817837012632e+17, 1.313817837034508e+17, 1.313817837057944e+17, 1.31381783707982e+17, 1.313817837103258e+17, 1.313817837125133e+17, 1.313817837147008e+17, 1.313817837170445e+17, 1.31381783719232e+17, 1.313817837215757e+17, 1.313817837237633e+17, 1.31381783726107e+17, 1.313817837282945e+17, 1.31381783730482e+17, 1.313817837328257e+17, 1.313817837350132e+17, 1.313817837381382e+17, 1.31381783740482e+17, 1.313817837428257e+17, 1.313817837450132e+17, 1.313817837473571e+17, 1.313817837495444e+17, 1.313817837518883e+17, 1.313817837540758e+17, 1.313817837562633e+17, 1.31381783758607e+17, 1.313817837607945e+17, 1.313817837631383e+17, 1.313817837653257e+17, 1.313817837676695e+17, 1.313817837707945e+17, 1.313817837731382e+17, 1.313817837753257e+17, 1.313817837776695e+17, 1.313817837798569e+17, 1.313817837820444e+17, 1.313817837843882e+17, 1.313817837865757e+17, 1.313817837889194e+17, 1.313817837911069e+17, 1.313817837934508e+17, 1.313817837956381e+17, 1.31381783797982e+17, 1.313817838001695e+17, 1.31381783802357e+17, 1.313817838047007e+17, 1.313817838068883e+17, 1.31381783809232e+17, 1.313817838115758e+17, 1.313817838147008e+17, 1.313817838168882e+17, 1.31381783819232e+17, 1.313817838215757e+17, 1.313817838237633e+17, 1.31381783826107e+17, 1.313817838282944e+17, 1.313817838306382e+17, 1.313817838328257e+17, 1.313817838350132e+17, 1.313817838373569e+17, 1.313817838395446e+17, 1.313817838418883e+17, 1.313817838440756e+17, 1.313817838473571e+17, 1.313817838495444e+17, 1.313817838518883e+17, 1.313817838540758e+17, 1.313817838564195e+17, 1.31381783858607e+17, 1.313817838607945e+17, 1.313817838631382e+17, 1.313817838653257e+17, 1.313817838676695e+17, 1.31381783869857e+17, 1.313817838722007e+17, 1.313817838743882e+17, 1.313817838765757e+17, 1.313817838789194e+17, 1.313817838811071e+17, 1.313817838834508e+17, 1.313817838856383e+17, 1.31381783887982e+17, 1.313817838911069e+17, 1.313817838934508e+17, 1.313817838956383e+17, 1.313817838979821e+17, 1.313817839003258e+17, 1.313817839025133e+17, 1.31381783904857e+17, 1.313817839072008e+17, 1.313817839093883e+17, 1.31381783911732e+17, 1.313817839140756e+17, 1.313817839162633e+17, 1.31381783918607e+17, 1.313817839209508e+17, 1.313817839239195e+17, 1.31381783926107e+17, 1.313817839284508e+17, 1.313817839306383e+17, 1.31381783932982e+17, 1.313817839351695e+17, 1.313817839375133e+17, 1.313817839397007e+17, 1.313817839418883e+17, 1.313817839442321e+17, 1.313817839464196e+17, 1.313817839487633e+17, 1.313817839509508e+17, 1.313817839532945e+17, 1.313817839562633e+17, 1.313817839584507e+17, 1.313817839607945e+17, 1.31381783962982e+17, 1.313817839653257e+17, 1.313817839676695e+17, 1.31381783969857e+17, 1.313817839722007e+17, 1.313817839743884e+17, 1.31381783976732e+17, 1.313817839789194e+17, 1.313817839811071e+17, 1.313817839834508e+17, 1.313817839856383e+17, 1.31381783987982e+17, 1.313817839903258e+17, 1.313817839925133e+17, 1.31381783994857e+17, 1.313817839970445e+17, 1.313817840003256e+17, 1.313817840026694e+17, 1.313817840050132e+17, 1.313817840072008e+17, 1.313817840095444e+17, 1.31381784011732e+17, 1.313817840140758e+17, 1.313817840162633e+17, 1.31381784018607e+17, 1.313817840207945e+17, 1.313817840231383e+17, 1.313817840253257e+17, 1.313817840275132e+17, 1.31381784029857e+17, 1.313817840331382e+17, 1.31381784035482e+17, 1.313817840376695e+17, 1.313817840398569e+17, 1.313817840422007e+17, 1.313817840443882e+17, 1.31381784046732e+17, 1.31381784049232e+17, 1.313817840514195e+17, 1.31381784053607e+17, 1.313817840559508e+17, 1.313817840581382e+17, 1.313817840604819e+17, 1.313817840628257e+17, 1.313817840657944e+17, 1.313817840681382e+17, 1.313817840703258e+17, 1.313817840725133e+17, 1.31381784074857e+17, 1.313817840770445e+17, 1.313817840793882e+17, 1.313817840815757e+17, 1.313817840839195e+17, 1.31381784086107e+17, 1.313817840884507e+17, 1.313817840906382e+17, 1.313817840928257e+17, 1.313817840951694e+17, 1.313817840981382e+17, 1.31381784100482e+17, 1.313817841028257e+17, 1.313817841050132e+17, 1.313817841073569e+17, 1.313817841097007e+17, 1.313817841118883e+17, 1.313817841142321e+17, 1.313817841164195e+17, 1.31381784118607e+17, 1.313817841209508e+17, 1.313817841232945e+17, 1.313817841256383e+17, 1.31381784127982e+17, 1.313817841312632e+17, 1.31381784133607e+17, 1.313817841359507e+17, 1.313817841382944e+17, 1.313817841406382e+17, 1.313817841428257e+17, 1.313817841451695e+17, 1.313817841475133e+17, 1.31381784149857e+17, 1.31381784152982e+17, 1.31381784155482e+17, 1.313817841578258e+17, 1.313817841601695e+17, 1.31381784162357e+17, 1.313817841647008e+17, 1.313817841672008e+17, 1.313817841693883e+17, 1.31381784171732e+17, 1.313817841750132e+17, 1.313817841772008e+17, 1.313817841795444e+17, 1.313817841817321e+17, 1.313817841839195e+17, 1.313817841862632e+17, 1.313817841884508e+17, 1.313817841907945e+17, 1.31381784192982e+17, 1.313817841953257e+17, 1.313817841975133e+17, 1.313817841997007e+17, 1.313817842020444e+17, 1.313817842042321e+17, 1.313817842065757e+17, 1.313817842087633e+17, 1.313817842111069e+17, 1.313817842132945e+17, 1.313817842156383e+17, 1.313817842187633e+17, 1.313817842211071e+17, 1.313817842232945e+17, 1.313817842256383e+17, 1.313817842278258e+17, 1.313817842300132e+17, 1.31381784232357e+17, 1.313817842345445e+17, 1.313817842368883e+17, 1.31381784239232e+17, 1.313817842414195e+17, 1.313817842437633e+17, 1.313817842459508e+17, 1.313817842482945e+17, 1.313817842514195e+17, 1.313817842537632e+17, 1.313817842559507e+17, 1.313817842581382e+17, 1.31381784260482e+17, 1.313817842626694e+17, 1.313817842650132e+17, 1.313817842672008e+17, 1.313817842695444e+17, 1.31381784271732e+17, 1.313817842740758e+17, 1.313817842762633e+17, 1.313817842784507e+17, 1.313817842807945e+17, 1.31381784282982e+17, 1.313817842853257e+17, 1.313817842875132e+17, 1.31381784289857e+17, 1.313817842920445e+17, 1.313817842951695e+17, 1.313817842973571e+17, 1.313817842997007e+17, 1.313817843018883e+17, 1.313817843042321e+17, 1.313817843065757e+17, 1.313817843090757e+17, 1.313817843115758e+17, 1.313817843181382e+17, 1.31381784320482e+17, 1.313817843226696e+17, 1.313817843250132e+17, 1.313817843272008e+17, 1.313817843295444e+17};
			mask_depths = {{15.0, 15.0, 51.6, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.4}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.4}, {15.0, 51.5}, {15.0, 51.4}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.4}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.5}, {15.0, 51.5}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.6}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.7}, {15.0, 51.7}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 52.0}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.8}, {15.0, 51.8}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.1}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.1}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.1}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 51.9}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 51.9}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.0}, {15.0, 51.9}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.0}, {15.0, 52.0}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.1}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.2}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.4}, {15.0, 52.3}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.3}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.3}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.3}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.4}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.5}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 15.0, 15.0, 15.0}};
		}
	}
}
