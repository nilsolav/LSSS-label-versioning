netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 14;
			channels = 4;
			categories = 56;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0, 81.1, 60.6, 65.7, 75.6, 68.9, 76.1, 75.9, 46.7, 71.2, 76.3, 76.3, 91.4, 60.0;
			max_depth =  93.9, 87.6, 65.4, 69.2, 78.4, 74.4, 80.2, 81.1, 51.6, 74.9, 91.3, 91.2, 93.9, 63.6;
			start_time = 129179007918085120, 129179012638710144, 129179010193241472, 129179008324491392, 129179010969022720, 129179014284022656, 129179013662460160, 129179014450585088, 129179012297460224, 129179015636835200, 129179019049335168, 129179019207772672, 129179019252460160, 129179007918085120;
			end_time = 129179019536991488, 129179012687460096, 129179010278397696, 129179008352772736, 129179010997460096, 129179014328710144, 129179013699022592, 129179014483085184, 129179012325897600, 129179015661210112, 129179019130585216, 129179019264647680, 129179019431210112, 129179007954647680;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14;
			region_name = "Layer1","Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "0", "0", "0", "0", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "0", "0", "0", "0", "27", "27", "27", "27";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "120", "200";
			region_channels = 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15;
			mask_times = {1.291790079180851e+17, 1.291790079221476e+17, 1.291790079262102e+17, 1.291790079302726e+17, 1.291790079343351e+17, 1.291790079383977e+17, 1.291790079424602e+17, 1.291790079465226e+17, 1.291790079505852e+17, 1.291790079546477e+17, 1.291790079587101e+17, 1.291790079627726e+17, 1.291790079668352e+17, 1.291790079708977e+17, 1.291790079749601e+17, 1.291790079790227e+17, 1.291790079830852e+17, 1.291790079871476e+17, 1.291790079912102e+17, 1.291790079952727e+17, 1.291790079993352e+17, 1.291790080033976e+17, 1.291790080074602e+17, 1.291790080115227e+17, 1.291790080155852e+17, 1.291790080196477e+17, 1.291790080237101e+17, 1.291790080277727e+17, 1.291790080318353e+17, 1.291790080358976e+17, 1.291790080399602e+17, 1.291790080440227e+17, 1.291790080480851e+17, 1.291790080521477e+17, 1.291790080562102e+17, 1.291790080602726e+17, 1.291790080643351e+17, 1.291790080683977e+17, 1.291790080724602e+17, 1.291790080765226e+17, 1.291790080805852e+17, 1.291790080846477e+17, 1.291790080887101e+17, 1.291790080927727e+17, 1.291790080968352e+17, 1.291790081008977e+17, 1.291790081049601e+17, 1.291790081090227e+17, 1.291790081130852e+17, 1.291790081171476e+17, 1.291790081212102e+17, 1.291790081252727e+17, 1.291790081293352e+17, 1.291790081333976e+17, 1.291790081374602e+17, 1.291790081415227e+17, 1.291790081455852e+17, 1.291790081496477e+17, 1.291790081537102e+17, 1.291790081577727e+17, 1.291790081616788e+17, 1.291790081658976e+17, 1.291790081699602e+17, 1.291790081740228e+17, 1.291790081780851e+17, 1.291790081821476e+17, 1.291790081862102e+17, 1.291790081902726e+17, 1.291790081943352e+17, 1.291790081983977e+17, 1.291790082026164e+17, 1.291790082066789e+17, 1.291790082107414e+17, 1.29179008214804e+17, 1.291790082188664e+17, 1.291790082227726e+17, 1.291790082269915e+17, 1.291790082308977e+17, 1.291790082351164e+17, 1.291790082390227e+17, 1.291790082432415e+17, 1.291790082473039e+17, 1.291790082513664e+17, 1.29179008255429e+17, 1.291790082594913e+17, 1.291790082635539e+17, 1.291790082676165e+17, 1.29179008271679e+17, 1.291790082757414e+17, 1.291790082798039e+17, 1.291790082838665e+17, 1.29179008287929e+17, 1.291790082919914e+17, 1.29179008296054e+17, 1.291790083001164e+17, 1.291790083041789e+17, 1.291790083080851e+17, 1.291790083121477e+17, 1.291790083162102e+17, 1.291790083204289e+17, 1.291790083244914e+17, 1.291790083283977e+17, 1.291790083324602e+17, 1.291790083365226e+17, 1.291790083405852e+17, 1.291790083446477e+17, 1.291790083487101e+17, 1.291790083527727e+17, 1.291790083568352e+17, 1.291790083608977e+17, 1.291790083649601e+17, 1.291790083690227e+17, 1.291790083730852e+17, 1.291790083773038e+17, 1.291790083813664e+17, 1.29179008385429e+17, 1.291790083893352e+17, 1.291790083933976e+17, 1.291790083974602e+17, 1.291790084015227e+17, 1.291790084055852e+17, 1.291790084096477e+17, 1.291790084137102e+17, 1.291790084177727e+17, 1.291790084218353e+17, 1.291790084258976e+17, 1.291790084299602e+17, 1.291790084340228e+17, 1.291790084380851e+17, 1.291790084421476e+17, 1.291790084462102e+17, 1.291790084505852e+17, 1.291790084546477e+17, 1.291790084587101e+17, 1.291790084627727e+17, 1.291790084668352e+17, 1.291790084707414e+17, 1.29179008474804e+17, 1.291790084788664e+17, 1.291790084829289e+17, 1.291790084869915e+17, 1.291790084912102e+17, 1.291790084951164e+17, 1.291790084991789e+17, 1.291790085032415e+17, 1.291790085073039e+17, 1.291790085113664e+17, 1.29179008515429e+17, 1.291790085194913e+17, 1.291790085235539e+17, 1.291790085277727e+17, 1.291790085316788e+17, 1.291790085358976e+17, 1.291790085398039e+17, 1.291790085438665e+17, 1.29179008547929e+17, 1.291790085519914e+17, 1.29179008556054e+17, 1.291790085601164e+17, 1.291790085641789e+17, 1.291790085682415e+17, 1.291790085723039e+17, 1.291790085763665e+17, 1.291790085804289e+17, 1.291790085844914e+17, 1.29179008588554e+17, 1.291790085926164e+17, 1.291790085966789e+17, 1.291790086007414e+17, 1.29179008604804e+17, 1.291790086088664e+17, 1.291790086127727e+17, 1.291790086168352e+17, 1.291790086208975e+17, 1.291790086249601e+17, 1.291790086290227e+17, 1.291790086330852e+17, 1.291790086371476e+17, 1.291790086412102e+17, 1.291790086452727e+17, 1.291790086493352e+17, 1.291790086533976e+17, 1.291790086577727e+17, 1.291790086616788e+17, 1.291790086657414e+17, 1.291790086698039e+17, 1.291790086738665e+17, 1.291790086779288e+17, 1.291790086819914e+17, 1.291790086858976e+17, 1.291790086899602e+17, 1.291790086940228e+17, 1.291790086980851e+17, 1.291790087021476e+17, 1.291790087062102e+17, 1.291790087102726e+17, 1.291790087143352e+17, 1.291790087183977e+17, 1.291790087224602e+17, 1.291790087265226e+17, 1.291790087305852e+17, 1.291790087346477e+17, 1.291790087387101e+17, 1.291790087427726e+17, 1.291790087468352e+17, 1.291790087508977e+17, 1.291790087549601e+17, 1.291790087590227e+17, 1.291790087630851e+17, 1.291790087671476e+17, 1.291790087712102e+17, 1.291790087752727e+17, 1.291790087793352e+17, 1.291790087833976e+17, 1.291790087874602e+17, 1.291790087915227e+17, 1.291790087955852e+17, 1.291790087996477e+17, 1.291790088037101e+17, 1.291790088077727e+17, 1.291790088118353e+17, 1.291790088158976e+17, 1.291790088199602e+17, 1.291790088240227e+17, 1.291790088280851e+17, 1.291790088321477e+17, 1.291790088362102e+17, 1.291790088402726e+17, 1.291790088441789e+17, 1.291790088483977e+17, 1.291790088524602e+17, 1.291790088565226e+17, 1.291790088605852e+17, 1.291790088646477e+17, 1.291790088687101e+17, 1.291790088727727e+17, 1.291790088768352e+17, 1.291790088808975e+17, 1.291790088849601e+17, 1.291790088890227e+17, 1.291790088930852e+17, 1.291790088971476e+17, 1.291790089012102e+17, 1.291790089052727e+17, 1.291790089093352e+17, 1.291790089133976e+17, 1.291790089174602e+17, 1.291790089215227e+17, 1.29179008925429e+17, 1.291790089296477e+17, 1.291790089337102e+17, 1.291790089377727e+17, 1.291790089418353e+17, 1.291790089458976e+17, 1.291790089499602e+17, 1.291790089540228e+17, 1.291790089580851e+17, 1.291790089621476e+17, 1.291790089662102e+17, 1.291790089702726e+17, 1.291790089743352e+17, 1.291790089783977e+17, 1.291790089824602e+17, 1.291790089865226e+17, 1.291790089905852e+17, 1.291790089946477e+17, 1.291790089987101e+17, 1.291790090027726e+17, 1.291790090068352e+17, 1.291790090108977e+17, 1.291790090149603e+17, 1.291790090190227e+17, 1.291790090230851e+17, 1.291790090271476e+17, 1.291790090312102e+17, 1.291790090352726e+17, 1.291790090393352e+17, 1.291790090433976e+17, 1.291790090474602e+17, 1.291790090515227e+17, 1.291790090555852e+17, 1.291790090596477e+17, 1.291790090637101e+17, 1.291790090677727e+17, 1.291790090716788e+17, 1.291790090758976e+17, 1.291790090799602e+17, 1.291790090840227e+17, 1.291790090880851e+17, 1.291790090919914e+17, 1.291790090960539e+17, 1.291790091002726e+17, 1.291790091043351e+17, 1.291790091083977e+17, 1.291790091124602e+17, 1.291790091165226e+17, 1.291790091205852e+17, 1.291790091246477e+17, 1.291790091287101e+17, 1.291790091327727e+17, 1.291790091368352e+17, 1.291790091408975e+17, 1.291790091449601e+17, 1.291790091490227e+17, 1.291790091530852e+17, 1.291790091571476e+17, 1.291790091612102e+17, 1.291790091652726e+17, 1.291790091693352e+17, 1.291790091733976e+17, 1.291790091774602e+17, 1.291790091815227e+17, 1.291790091855852e+17, 1.291790091896477e+17, 1.291790091937102e+17, 1.291790091977727e+17, 1.291790092018353e+17, 1.291790092058976e+17, 1.291790092099602e+17, 1.291790092140228e+17, 1.291790092180851e+17, 1.291790092221476e+17, 1.291790092262102e+17, 1.291790092302726e+17, 1.291790092343352e+17, 1.291790092383977e+17, 1.291790092424602e+17, 1.291790092465226e+17, 1.291790092505852e+17, 1.291790092546477e+17, 1.291790092587101e+17, 1.291790092627726e+17, 1.291790092668352e+17, 1.291790092708977e+17, 1.291790092749603e+17, 1.291790092790227e+17, 1.291790092830851e+17, 1.291790092871476e+17, 1.291790092912102e+17, 1.291790092952726e+17, 1.291790092993352e+17, 1.291790093033976e+17, 1.291790093074601e+17, 1.291790093115227e+17, 1.291790093155852e+17, 1.291790093196477e+17, 1.291790093237101e+17, 1.291790093277727e+17, 1.291790093318353e+17, 1.291790093358976e+17, 1.291790093399602e+17, 1.291790093440227e+17, 1.291790093480851e+17, 1.291790093521477e+17, 1.291790093562102e+17, 1.291790093602726e+17, 1.291790093643351e+17, 1.291790093683977e+17, 1.291790093724602e+17, 1.291790093765226e+17, 1.291790093805852e+17, 1.291790093846477e+17, 1.291790093887101e+17, 1.291790093927727e+17, 1.291790093968352e+17, 1.291790094008977e+17, 1.291790094049601e+17, 1.291790094090227e+17, 1.291790094129289e+17, 1.291790094171476e+17, 1.291790094212102e+17, 1.291790094252726e+17, 1.291790094293352e+17, 1.291790094333978e+17, 1.291790094374601e+17, 1.291790094415227e+17, 1.291790094455852e+17, 1.291790094496476e+17, 1.291790094537102e+17, 1.291790094577727e+17, 1.291790094618353e+17, 1.291790094658976e+17, 1.291790094699602e+17, 1.291790094740228e+17, 1.291790094780851e+17, 1.291790094821476e+17, 1.291790094862102e+17, 1.291790094902726e+17, 1.291790094943352e+17, 1.291790094983977e+17, 1.291790095024602e+17, 1.291790095065226e+17, 1.291790095105852e+17, 1.291790095146477e+17, 1.291790095187101e+17, 1.291790095227727e+17, 1.291790095268352e+17, 1.291790095308977e+17, 1.291790095349603e+17, 1.291790095390227e+17, 1.291790095430851e+17, 1.291790095471476e+17, 1.291790095512102e+17, 1.291790095552727e+17, 1.291790095593352e+17, 1.291790095633976e+17, 1.291790095674601e+17, 1.291790095715227e+17, 1.291790095755852e+17, 1.291790095796476e+17, 1.291790095837101e+17, 1.291790095877727e+17, 1.291790095918353e+17, 1.291790095958976e+17, 1.291790095999602e+17, 1.291790096040227e+17, 1.291790096080851e+17, 1.291790096121477e+17, 1.291790096162102e+17, 1.291790096202726e+17, 1.291790096243351e+17, 1.291790096283977e+17, 1.291790096326164e+17, 1.291790096366789e+17, 1.291790096405852e+17, 1.291790096446477e+17, 1.291790096487101e+17, 1.291790096527727e+17, 1.291790096568352e+17, 1.291790096608977e+17, 1.291790096649601e+17, 1.291790096690227e+17, 1.291790096730852e+17, 1.291790096771476e+17, 1.291790096812102e+17, 1.291790096852726e+17, 1.291790096893352e+17, 1.291790096933978e+17, 1.291790096974601e+17, 1.291790097015227e+17, 1.291790097055852e+17, 1.291790097096476e+17, 1.291790097137102e+17, 1.291790097177727e+17, 1.291790097216788e+17, 1.291790097258976e+17, 1.291790097299602e+17, 1.291790097340228e+17, 1.291790097380851e+17, 1.291790097421476e+17, 1.291790097462102e+17, 1.291790097502726e+17, 1.291790097543352e+17, 1.291790097583977e+17, 1.291790097624602e+17, 1.291790097665226e+17, 1.291790097705852e+17, 1.29179009774804e+17, 1.291790097787101e+17, 1.291790097827727e+17, 1.291790097868352e+17, 1.291790097908977e+17, 1.291790097949603e+17, 1.291790097990227e+17, 1.291790098030852e+17, 1.291790098071476e+17, 1.291790098112102e+17, 1.291790098152727e+17, 1.291790098193352e+17, 1.291790098233976e+17, 1.291790098274601e+17, 1.291790098315227e+17, 1.291790098355853e+17, 1.291790098396476e+17, 1.291790098437101e+17, 1.291790098477727e+17, 1.291790098518351e+17, 1.291790098558976e+17, 1.291790098599602e+17, 1.291790098640227e+17, 1.29179009867929e+17, 1.291790098721477e+17, 1.291790098762102e+17, 1.291790098802726e+17, 1.291790098843351e+17, 1.291790098883977e+17, 1.291790098924602e+17, 1.291790098965226e+17, 1.291790099005852e+17, 1.291790099046477e+17, 1.291790099087101e+17, 1.291790099127727e+17, 1.291790099168352e+17, 1.291790099208977e+17, 1.291790099249601e+17, 1.291790099290227e+17, 1.291790099330852e+17, 1.291790099371476e+17, 1.291790099412102e+17, 1.291790099452726e+17, 1.291790099493352e+17, 1.291790099533978e+17, 1.291790099574601e+17, 1.291790099615227e+17, 1.291790099655852e+17, 1.291790099696476e+17, 1.291790099737102e+17, 1.291790099777727e+17, 1.291790099818351e+17, 1.291790099858976e+17, 1.291790099899602e+17, 1.291790099940227e+17, 1.291790099980851e+17, 1.291790100021476e+17, 1.291790100062102e+17, 1.291790100102726e+17, 1.291790100143352e+17, 1.291790100183977e+17, 1.291790100224602e+17, 1.291790100265226e+17, 1.291790100305852e+17, 1.291790100346477e+17, 1.291790100387101e+17, 1.291790100427727e+17, 1.291790100468352e+17, 1.291790100508977e+17, 1.291790100549603e+17, 1.291790100590227e+17, 1.291790100629289e+17, 1.291790100671476e+17, 1.291790100712102e+17, 1.291790100752727e+17, 1.291790100793352e+17, 1.291790100833976e+17, 1.291790100874601e+17, 1.291790100915227e+17, 1.291790100955853e+17, 1.291790100996476e+17, 1.291790101037101e+17, 1.291790101077727e+17, 1.291790101118351e+17, 1.291790101158976e+17, 1.291790101199602e+17, 1.291790101240227e+17, 1.291790101280851e+17, 1.291790101321477e+17, 1.291790101362102e+17, 1.291790101402726e+17, 1.291790101443351e+17, 1.291790101483977e+17, 1.291790101524602e+17, 1.291790101565226e+17, 1.291790101605852e+17, 1.291790101646477e+17, 1.291790101687101e+17, 1.291790101727727e+17, 1.291790101768352e+17, 1.291790101808977e+17, 1.291790101851164e+17, 1.291790101890227e+17, 1.291790101932415e+17, 1.291790101971476e+17, 1.291790102012102e+17, 1.291790102052726e+17, 1.291790102093352e+17, 1.291790102133978e+17, 1.291790102174601e+17, 1.291790102215227e+17, 1.291790102255852e+17, 1.291790102296476e+17, 1.291790102337102e+17, 1.291790102377727e+17, 1.291790102418351e+17, 1.291790102458976e+17, 1.291790102499602e+17, 1.291790102540227e+17, 1.291790102580851e+17, 1.291790102621476e+17, 1.291790102662102e+17, 1.291790102702726e+17, 1.291790102743352e+17, 1.291790102783977e+17, 1.291790102824602e+17, 1.291790102865226e+17, 1.291790102905852e+17, 1.291790102946477e+17, 1.291790102987101e+17, 1.291790103027727e+17, 1.291790103068352e+17, 1.291790103108977e+17, 1.291790103149603e+17, 1.291790103190227e+17, 1.291790103230852e+17, 1.291790103271476e+17, 1.291790103312102e+17, 1.291790103352727e+17, 1.291790103393352e+17, 1.291790103433976e+17, 1.291790103474601e+17, 1.291790103515227e+17, 1.291790103555853e+17, 1.291790103596476e+17, 1.291790103637101e+17, 1.291790103677727e+17, 1.291790103718351e+17, 1.291790103758976e+17, 1.291790103799602e+17, 1.291790103840227e+17, 1.291790103880851e+17, 1.291790103921477e+17, 1.291790103962102e+17, 1.291790104002726e+17, 1.291790104041789e+17, 1.291790104083977e+17, 1.291790104124602e+17, 1.291790104165226e+17, 1.291790104205852e+17, 1.291790104246477e+17, 1.291790104287101e+17, 1.291790104327727e+17, 1.291790104369915e+17, 1.291790104408977e+17, 1.291790104449601e+17, 1.291790104490227e+17, 1.291790104530852e+17, 1.291790104571476e+17, 1.291790104612102e+17, 1.291790104652726e+17, 1.291790104693352e+17, 1.291790104733978e+17, 1.291790104774601e+17, 1.291790104815227e+17, 1.291790104855852e+17, 1.291790104896476e+17, 1.291790104937102e+17, 1.291790104977727e+17, 1.291790105018351e+17, 1.291790105058976e+17, 1.291790105099602e+17, 1.291790105140227e+17, 1.291790105180851e+17, 1.291790105221476e+17, 1.291790105262102e+17, 1.291790105302726e+17, 1.291790105343352e+17, 1.291790105383977e+17, 1.291790105424602e+17, 1.291790105465226e+17, 1.291790105505852e+17, 1.291790105546477e+17, 1.291790105587101e+17, 1.291790105627727e+17, 1.291790105668352e+17, 1.291790105708977e+17, 1.291790105749603e+17, 1.291790105790227e+17, 1.291790105830852e+17, 1.291790105871476e+17, 1.291790105912102e+17, 1.291790105952727e+17, 1.291790105993352e+17, 1.291790106033976e+17, 1.291790106074601e+17, 1.291790106115227e+17, 1.291790106155853e+17, 1.291790106196476e+17, 1.291790106237102e+17, 1.291790106277727e+17, 1.291790106318351e+17, 1.291790106358976e+17, 1.291790106399602e+17, 1.291790106440227e+17, 1.291790106480851e+17, 1.291790106521477e+17, 1.291790106562102e+17, 1.291790106602726e+17, 1.291790106641789e+17, 1.291790106683977e+17, 1.291790106724602e+17, 1.291790106765226e+17, 1.291790106805852e+17, 1.291790106846477e+17, 1.291790106887101e+17, 1.291790106927727e+17, 1.291790106968352e+17, 1.291790107008977e+17, 1.291790107049601e+17, 1.291790107090227e+17, 1.291790107130852e+17, 1.291790107171476e+17, 1.291790107212102e+17, 1.291790107252726e+17, 1.291790107293352e+17, 1.291790107333978e+17, 1.291790107374601e+17, 1.291790107415227e+17, 1.291790107455852e+17, 1.291790107496476e+17, 1.291790107537102e+17, 1.291790107577727e+17, 1.291790107618351e+17, 1.291790107658976e+17, 1.291790107699602e+17, 1.291790107740227e+17, 1.291790107780851e+17, 1.291790107821476e+17, 1.291790107862102e+17, 1.291790107902726e+17, 1.291790107943352e+17, 1.291790107983977e+17, 1.291790108024602e+17, 1.291790108065226e+17, 1.291790108105852e+17, 1.291790108146477e+17, 1.291790108187101e+17, 1.291790108227727e+17, 1.291790108268352e+17, 1.291790108308977e+17, 1.291790108349603e+17, 1.291790108390227e+17, 1.291790108430852e+17, 1.291790108471476e+17, 1.291790108512102e+17, 1.291790108552727e+17, 1.291790108593352e+17, 1.291790108633976e+17, 1.291790108674601e+17, 1.291790108715227e+17, 1.291790108755853e+17, 1.291790108796476e+17, 1.291790108837102e+17, 1.291790108877727e+17, 1.291790108918351e+17, 1.291790108958976e+17, 1.291790108999602e+17, 1.291790109040227e+17, 1.291790109080851e+17, 1.291790109121477e+17, 1.291790109162102e+17, 1.291790109202726e+17, 1.291790109243351e+17, 1.291790109283977e+17, 1.291790109324602e+17, 1.291790109365228e+17, 1.291790109405852e+17, 1.291790109446477e+17, 1.291790109487101e+17, 1.291790109527727e+17, 1.291790109568352e+17, 1.291790109608977e+17, 1.291790109649601e+17, 1.291790109690227e+17, 1.291790109729289e+17, 1.291790109769915e+17, 1.291790109812102e+17, 1.291790109852726e+17, 1.291790109893352e+17, 1.291790109933978e+17, 1.291790109974601e+17, 1.291790110015227e+17, 1.291790110055852e+17, 1.291790110096476e+17, 1.291790110137102e+17, 1.291790110177727e+17, 1.291790110218351e+17, 1.291790110258976e+17, 1.291790110299602e+17, 1.291790110340227e+17, 1.291790110380851e+17, 1.291790110421477e+17, 1.291790110462102e+17, 1.291790110502726e+17, 1.291790110543352e+17, 1.291790110583977e+17, 1.291790110624602e+17, 1.291790110665226e+17, 1.291790110705852e+17, 1.291790110746477e+17, 1.291790110787101e+17, 1.291790110827727e+17, 1.291790110868352e+17, 1.291790110908977e+17, 1.291790110949603e+17, 1.291790110990227e+17, 1.291790111030852e+17, 1.291790111071476e+17, 1.291790111112102e+17, 1.291790111152727e+17, 1.291790111193352e+17, 1.291790111233976e+17, 1.291790111274601e+17, 1.291790111315227e+17, 1.291790111355853e+17, 1.291790111396476e+17, 1.291790111437102e+17, 1.291790111477727e+17, 1.291790111518351e+17, 1.291790111558976e+17, 1.291790111599602e+17, 1.291790111640227e+17, 1.291790111680851e+17, 1.291790111721477e+17, 1.291790111762102e+17, 1.291790111802726e+17, 1.291790111843351e+17, 1.291790111883977e+17, 1.291790111924602e+17, 1.291790111965228e+17, 1.291790112005852e+17, 1.291790112044914e+17, 1.291790112087101e+17, 1.291790112127727e+17, 1.291790112168352e+17, 1.291790112208977e+17, 1.291790112249601e+17, 1.291790112290227e+17, 1.291790112330852e+17, 1.291790112371476e+17, 1.291790112412102e+17, 1.291790112452726e+17, 1.291790112493352e+17, 1.291790112533978e+17, 1.291790112574601e+17, 1.291790112615227e+17, 1.291790112655852e+17, 1.291790112696476e+17, 1.291790112737102e+17, 1.291790112777727e+17, 1.291790112818351e+17, 1.291790112858976e+17, 1.291790112899602e+17, 1.291790112940227e+17, 1.291790112980851e+17, 1.291790113021477e+17, 1.291790113062102e+17, 1.291790113102726e+17, 1.291790113141789e+17, 1.291790113183977e+17, 1.291790113224602e+17, 1.291790113265226e+17, 1.291790113305852e+17, 1.291790113346477e+17, 1.291790113387101e+17, 1.291790113427727e+17, 1.291790113468352e+17, 1.291790113508977e+17, 1.291790113549603e+17, 1.291790113590227e+17, 1.291790113630852e+17, 1.291790113671476e+17, 1.291790113712102e+17, 1.291790113752727e+17, 1.291790113793352e+17, 1.291790113833976e+17, 1.291790113874601e+17, 1.291790113915227e+17, 1.291790113955853e+17, 1.291790113996476e+17, 1.291790114037102e+17, 1.291790114077727e+17, 1.291790114118351e+17, 1.291790114158976e+17, 1.291790114199602e+17, 1.291790114240227e+17, 1.291790114280851e+17, 1.291790114321477e+17, 1.291790114362102e+17, 1.291790114402726e+17, 1.291790114443352e+17, 1.291790114483977e+17, 1.291790114524602e+17, 1.291790114565228e+17, 1.291790114605852e+17, 1.291790114646476e+17, 1.291790114687101e+17, 1.291790114727727e+17, 1.291790114768352e+17, 1.291790114808977e+17, 1.29179011484804e+17, 1.291790114890227e+17, 1.291790114930852e+17, 1.291790114973039e+17, 1.291790115012102e+17, 1.291790115052726e+17, 1.291790115093352e+17, 1.291790115133978e+17, 1.291790115174601e+17, 1.291790115215227e+17, 1.291790115255852e+17, 1.291790115296476e+17, 1.291790115337102e+17, 1.291790115377727e+17, 1.291790115416788e+17, 1.291790115458976e+17, 1.291790115499602e+17, 1.291790115540227e+17, 1.291790115580851e+17, 1.291790115621477e+17, 1.291790115662102e+17, 1.291790115702726e+17, 1.291790115741789e+17, 1.291790115783977e+17, 1.291790115824602e+17, 1.291790115865226e+17, 1.291790115905852e+17, 1.291790115946477e+17, 1.291790115987101e+17, 1.291790116027727e+17, 1.291790116068351e+17, 1.291790116108977e+17, 1.291790116149603e+17, 1.291790116190227e+17, 1.291790116230852e+17, 1.291790116271476e+17, 1.291790116312102e+17, 1.291790116352727e+17, 1.291790116393352e+17, 1.291790116433976e+17, 1.291790116474601e+17, 1.291790116515227e+17, 1.291790116555853e+17, 1.291790116596476e+17, 1.291790116637102e+17, 1.291790116677727e+17, 1.291790116718351e+17, 1.291790116758976e+17, 1.291790116799602e+17, 1.291790116840227e+17, 1.291790116880851e+17, 1.291790116921477e+17, 1.291790116962102e+17, 1.291790117002726e+17, 1.291790117043352e+17, 1.291790117083977e+17, 1.291790117124602e+17, 1.291790117165228e+17, 1.291790117205852e+17, 1.291790117246476e+17, 1.291790117287101e+17, 1.291790117327727e+17, 1.291790117368352e+17, 1.291790117408977e+17, 1.291790117449601e+17, 1.291790117490226e+17, 1.291790117530852e+17, 1.291790117571476e+17, 1.291790117612102e+17, 1.291790117652726e+17, 1.291790117693352e+17, 1.291790117733978e+17, 1.291790117774601e+17, 1.291790117815227e+17, 1.291790117855852e+17, 1.291790117896476e+17, 1.291790117937102e+17, 1.291790117977727e+17, 1.291790118016788e+17, 1.291790118058976e+17, 1.291790118099602e+17, 1.291790118140227e+17, 1.291790118180851e+17, 1.291790118221477e+17, 1.291790118262102e+17, 1.291790118302726e+17, 1.291790118343352e+17, 1.291790118383977e+17, 1.291790118424602e+17, 1.291790118465226e+17, 1.291790118505852e+17, 1.291790118546477e+17, 1.291790118587101e+17, 1.291790118627727e+17, 1.291790118668351e+17, 1.291790118708977e+17, 1.291790118749603e+17, 1.291790118790226e+17, 1.291790118830852e+17, 1.291790118871476e+17, 1.291790118912102e+17, 1.291790118952727e+17, 1.291790118993352e+17, 1.291790119033976e+17, 1.291790119074601e+17, 1.291790119115227e+17, 1.291790119155853e+17, 1.291790119196476e+17, 1.291790119237102e+17, 1.291790119277727e+17, 1.291790119318351e+17, 1.291790119358976e+17, 1.291790119399602e+17, 1.291790119440227e+17, 1.291790119480851e+17, 1.291790119521477e+17, 1.291790119562102e+17, 1.291790119602726e+17, 1.291790119643352e+17, 1.291790119683977e+17, 1.291790119724602e+17, 1.291790119765228e+17, 1.291790119805852e+17, 1.291790119846476e+17, 1.291790119887101e+17, 1.291790119927727e+17, 1.291790119968352e+17, 1.291790120008977e+17, 1.291790120049601e+17, 1.291790120090226e+17, 1.291790120130852e+17, 1.291790120171476e+17, 1.291790120212101e+17, 1.291790120252726e+17, 1.291790120291789e+17, 1.291790120333978e+17, 1.291790120374601e+17, 1.291790120415227e+17, 1.291790120455852e+17, 1.291790120496476e+17, 1.291790120537102e+17, 1.291790120577727e+17, 1.291790120618351e+17, 1.291790120658976e+17, 1.291790120699602e+17, 1.291790120740227e+17, 1.291790120780851e+17, 1.291790120821477e+17, 1.291790120862102e+17, 1.291790120902726e+17, 1.291790120943352e+17, 1.291790120983977e+17, 1.291790121024602e+17, 1.291790121065226e+17, 1.291790121105852e+17, 1.291790121144914e+17, 1.291790121187101e+17, 1.291790121227727e+17, 1.291790121268351e+17, 1.291790121308977e+17, 1.291790121349603e+17, 1.291790121390226e+17, 1.291790121429289e+17, 1.291790121471476e+17, 1.291790121512101e+17, 1.291790121552727e+17, 1.291790121593352e+17, 1.291790121633976e+17, 1.291790121674601e+17, 1.291790121715227e+17, 1.291790121755853e+17, 1.291790121796476e+17, 1.291790121837102e+17, 1.291790121877727e+17, 1.291790121918351e+17, 1.291790121958976e+17, 1.291790121999602e+17, 1.291790122040227e+17, 1.291790122080851e+17, 1.291790122121477e+17, 1.291790122162102e+17, 1.291790122202726e+17, 1.291790122243352e+17, 1.291790122283977e+17, 1.291790122324602e+17, 1.291790122365228e+17, 1.291790122405852e+17, 1.291790122446476e+17, 1.291790122487101e+17, 1.291790122527727e+17, 1.291790122568352e+17, 1.291790122608977e+17, 1.291790122649603e+17, 1.291790122690226e+17, 1.291790122730852e+17, 1.291790122771476e+17, 1.291790122812101e+17, 1.291790122852726e+17, 1.291790122893352e+17, 1.291790122933976e+17, 1.291790122974602e+17, 1.291790123015227e+17, 1.291790123055852e+17, 1.291790123096476e+17, 1.291790123137102e+17, 1.291790123177727e+17, 1.291790123218351e+17, 1.291790123258976e+17, 1.291790123299602e+17, 1.291790123340227e+17, 1.291790123380851e+17, 1.291790123421477e+17, 1.291790123462102e+17, 1.291790123502726e+17, 1.291790123543352e+17, 1.291790123583977e+17, 1.291790123624602e+17, 1.291790123665226e+17, 1.291790123705852e+17, 1.291790123746477e+17, 1.291790123787101e+17, 1.291790123827727e+17, 1.291790123868351e+17, 1.291790123908977e+17, 1.291790123949603e+17, 1.291790123990226e+17, 1.291790124030852e+17, 1.291790124073039e+17, 1.291790124112101e+17, 1.291790124152727e+17, 1.291790124193352e+17, 1.291790124233976e+17, 1.291790124274601e+17, 1.291790124315227e+17, 1.291790124355852e+17, 1.291790124396476e+17, 1.291790124437102e+17, 1.291790124477727e+17, 1.291790124518351e+17, 1.291790124558976e+17, 1.291790124599602e+17, 1.291790124640227e+17, 1.291790124680851e+17, 1.291790124721477e+17, 1.291790124762102e+17, 1.291790124802726e+17, 1.291790124843352e+17, 1.291790124883977e+17, 1.291790124924602e+17, 1.291790124965228e+17, 1.291790125005852e+17, 1.291790125046476e+17, 1.291790125087101e+17, 1.291790125127727e+17, 1.291790125168352e+17, 1.291790125208977e+17, 1.291790125249603e+17, 1.291790125290226e+17, 1.291790125330852e+17, 1.291790125371476e+17, 1.291790125412101e+17, 1.291790125452727e+17, 1.291790125493352e+17, 1.291790125533976e+17, 1.291790125574602e+17, 1.291790125615227e+17, 1.291790125655852e+17, 1.291790125698039e+17, 1.291790125737102e+17, 1.291790125777728e+17, 1.291790125818351e+17, 1.291790125858976e+17, 1.291790125899602e+17, 1.291790125940227e+17, 1.29179012597929e+17, 1.291790126023039e+17, 1.291790126062102e+17, 1.291790126102726e+17, 1.291790126143352e+17, 1.291790126183977e+17, 1.291790126224602e+17, 1.291790126265226e+17, 1.291790126305852e+17, 1.291790126346477e+17, 1.291790126387101e+17, 1.291790126427727e+17, 1.291790126468351e+17, 1.291790126508977e+17, 1.291790126549603e+17, 1.291790126590226e+17, 1.291790126630852e+17, 1.291790126671476e+17, 1.291790126712101e+17, 1.291790126752727e+17, 1.291790126793352e+17, 1.291790126833976e+17, 1.291790126874601e+17, 1.291790126915227e+17, 1.291790126955852e+17, 1.291790126996476e+17, 1.291790127037102e+17, 1.291790127077727e+17, 1.291790127118351e+17, 1.291790127158977e+17, 1.291790127199602e+17, 1.291790127240227e+17, 1.291790127280851e+17, 1.291790127321477e+17, 1.291790127362102e+17, 1.291790127402726e+17, 1.291790127443352e+17, 1.291790127483977e+17, 1.291790127526164e+17, 1.291790127565228e+17, 1.291790127605852e+17, 1.291790127646476e+17, 1.291790127687101e+17, 1.291790127727727e+17, 1.291790127768352e+17, 1.291790127808977e+17, 1.291790127849603e+17, 1.291790127890226e+17, 1.291790127930852e+17, 1.291790127971476e+17, 1.291790128012101e+17, 1.291790128052727e+17, 1.291790128093352e+17, 1.291790128133976e+17, 1.291790128174602e+17, 1.291790128215227e+17, 1.291790128255852e+17, 1.291790128296476e+17, 1.291790128337102e+17, 1.291790128377727e+17, 1.291790128418351e+17, 1.291790128458976e+17, 1.291790128499602e+17, 1.291790128540227e+17, 1.291790128580851e+17, 1.291790128621477e+17, 1.291790128662102e+17, 1.291790128702726e+17, 1.291790128743352e+17, 1.291790128783977e+17, 1.291790128824602e+17, 1.291790128865226e+17, 1.291790128905852e+17, 1.291790128946477e+17, 1.291790128987101e+17, 1.291790129027727e+17, 1.291790129068351e+17, 1.291790129108977e+17, 1.291790129149603e+17, 1.291790129190226e+17, 1.291790129230852e+17, 1.291790129271476e+17, 1.291790129312101e+17, 1.291790129352727e+17, 1.291790129393352e+17, 1.291790129433976e+17, 1.291790129474601e+17, 1.291790129515227e+17, 1.291790129555852e+17, 1.291790129596476e+17, 1.291790129637102e+17, 1.291790129677727e+17, 1.291790129718351e+17, 1.291790129758977e+17, 1.291790129799602e+17, 1.291790129840227e+17, 1.291790129880851e+17, 1.291790129921477e+17, 1.291790129962102e+17, 1.291790130002726e+17, 1.291790130044914e+17, 1.29179013008554e+17, 1.291790130124602e+17, 1.291790130165228e+17, 1.291790130205852e+17, 1.291790130246476e+17, 1.291790130287101e+17, 1.291790130327727e+17, 1.291790130368352e+17, 1.291790130408977e+17, 1.291790130449603e+17, 1.291790130490226e+17, 1.291790130530852e+17, 1.291790130571476e+17, 1.291790130612101e+17, 1.291790130652727e+17, 1.291790130693352e+17, 1.291790130733976e+17, 1.291790130774602e+17, 1.291790130815227e+17, 1.291790130855852e+17, 1.291790130896476e+17, 1.291790130937102e+17, 1.291790130977727e+17, 1.291790131018351e+17, 1.291790131058976e+17, 1.291790131099602e+17, 1.291790131140227e+17, 1.291790131180852e+17, 1.291790131221477e+17, 1.291790131262102e+17, 1.291790131302726e+17, 1.291790131343352e+17, 1.291790131383977e+17, 1.291790131424602e+17, 1.291790131465226e+17, 1.291790131505852e+17, 1.291790131546477e+17, 1.291790131587101e+17, 1.291790131627727e+17, 1.291790131668351e+17, 1.291790131708977e+17, 1.291790131749603e+17, 1.291790131790226e+17, 1.291790131830852e+17, 1.291790131871476e+17, 1.291790131912101e+17, 1.291790131952727e+17, 1.291790131993352e+17, 1.291790132035539e+17, 1.291790132074601e+17, 1.291790132115227e+17, 1.291790132155852e+17, 1.291790132196476e+17, 1.291790132237102e+17, 1.291790132277727e+17, 1.291790132318351e+17, 1.291790132358977e+17, 1.291790132399602e+17, 1.291790132440227e+17, 1.291790132480851e+17, 1.291790132521477e+17, 1.291790132562102e+17, 1.291790132602726e+17, 1.291790132643352e+17, 1.291790132683977e+17, 1.291790132724602e+17, 1.291790132765228e+17, 1.291790132805852e+17, 1.291790132846476e+17, 1.291790132887101e+17, 1.291790132927727e+17, 1.291790132968352e+17, 1.291790133008977e+17, 1.291790133049603e+17, 1.291790133090226e+17, 1.291790133132413e+17, 1.291790133171476e+17, 1.291790133212101e+17, 1.291790133252727e+17, 1.291790133293352e+17, 1.291790133333976e+17, 1.291790133374602e+17, 1.291790133415227e+17, 1.291790133455852e+17, 1.291790133496476e+17, 1.291790133537102e+17, 1.291790133577727e+17, 1.291790133618351e+17, 1.291790133658976e+17, 1.291790133699602e+17, 1.291790133740227e+17, 1.291790133780852e+17, 1.291790133821477e+17, 1.291790133862102e+17, 1.291790133902726e+17, 1.291790133943352e+17, 1.291790133983977e+17, 1.291790134024602e+17, 1.291790134065226e+17, 1.291790134105852e+17, 1.291790134146477e+17, 1.29179013418554e+17, 1.291790134227727e+17, 1.291790134268351e+17, 1.291790134308977e+17, 1.291790134349603e+17, 1.291790134390226e+17, 1.291790134430852e+17, 1.291790134471476e+17, 1.291790134512101e+17, 1.291790134552727e+17, 1.291790134593352e+17, 1.291790134633976e+17, 1.291790134674601e+17, 1.291790134715227e+17, 1.291790134755852e+17, 1.291790134796476e+17, 1.291790134837102e+17, 1.291790134877727e+17, 1.291790134918351e+17, 1.291790134958977e+17, 1.291790134999602e+17, 1.291790135040227e+17, 1.29179013507929e+17, 1.291790135121477e+17, 1.291790135162102e+17, 1.291790135202726e+17, 1.291790135243352e+17, 1.291790135283977e+17, 1.291790135324602e+17, 1.291790135365228e+17, 1.291790135405852e+17, 1.291790135446476e+17, 1.291790135487101e+17, 1.291790135527727e+17, 1.291790135568352e+17, 1.291790135608977e+17, 1.291790135649603e+17, 1.291790135690226e+17, 1.291790135730852e+17, 1.291790135771476e+17, 1.291790135812101e+17, 1.291790135852727e+17, 1.291790135891789e+17, 1.291790135933976e+17, 1.291790135974602e+17, 1.291790136015227e+17, 1.291790136055852e+17, 1.291790136096476e+17, 1.291790136137102e+17, 1.291790136177727e+17, 1.29179013621679e+17, 1.291790136258976e+17, 1.291790136299602e+17, 1.291790136340227e+17, 1.291790136380852e+17, 1.291790136421477e+17, 1.291790136462102e+17, 1.291790136502726e+17, 1.291790136543352e+17, 1.291790136583977e+17, 1.291790136624602e+17, 1.291790136665226e+17, 1.291790136705852e+17, 1.291790136746477e+17, 1.291790136787103e+17, 1.291790136827727e+17, 1.291790136868351e+17, 1.291790136908977e+17, 1.291790136949603e+17, 1.291790136990226e+17, 1.29179013702929e+17, 1.291790137071476e+17, 1.291790137112101e+17, 1.291790137152727e+17, 1.291790137193352e+17, 1.291790137233976e+17, 1.291790137274601e+17, 1.291790137315227e+17, 1.291790137355852e+17, 1.291790137396476e+17, 1.291790137437102e+17, 1.291790137477727e+17, 1.291790137518351e+17, 1.291790137558977e+17, 1.291790137599602e+17, 1.291790137640227e+17, 1.291790137680851e+17, 1.291790137721477e+17, 1.291790137762102e+17, 1.291790137802726e+17, 1.291790137843352e+17, 1.291790137883977e+17, 1.291790137924602e+17, 1.291790137965228e+17, 1.291790138005852e+17, 1.291790138046476e+17, 1.291790138087101e+17, 1.291790138127727e+17, 1.291790138168352e+17, 1.291790138208977e+17, 1.291790138249603e+17, 1.291790138290226e+17, 1.291790138330852e+17, 1.291790138371476e+17, 1.291790138412101e+17, 1.291790138452727e+17, 1.291790138491789e+17, 1.291790138533976e+17, 1.291790138574602e+17, 1.291790138615227e+17, 1.291790138655852e+17, 1.291790138696476e+17, 1.291790138737102e+17, 1.291790138777727e+17, 1.291790138818351e+17, 1.291790138858976e+17, 1.291790138899602e+17, 1.291790138940227e+17, 1.291790138980852e+17, 1.291790139021477e+17, 1.291790139062102e+17, 1.291790139102726e+17, 1.291790139143352e+17, 1.291790139183976e+17, 1.291790139224602e+17, 1.291790139265226e+17, 1.291790139305852e+17, 1.291790139344914e+17, 1.291790139387103e+17, 1.291790139427727e+17, 1.291790139468351e+17, 1.291790139508977e+17, 1.291790139549603e+17, 1.291790139590226e+17, 1.291790139630852e+17, 1.291790139671476e+17, 1.291790139712101e+17, 1.291790139752727e+17, 1.291790139793352e+17, 1.291790139833976e+17, 1.291790139874601e+17, 1.291790139915227e+17, 1.291790139955852e+17, 1.291790139996476e+17, 1.291790140037102e+17, 1.291790140077727e+17, 1.291790140118351e+17, 1.291790140158977e+17, 1.291790140199602e+17, 1.291790140240227e+17, 1.291790140280851e+17, 1.291790140321477e+17, 1.291790140362102e+17, 1.291790140402726e+17, 1.291790140443352e+17, 1.291790140483976e+17, 1.291790140524602e+17, 1.291790140565228e+17, 1.291790140605852e+17, 1.291790140648038e+17, 1.291790140687101e+17, 1.291790140727727e+17, 1.291790140768352e+17, 1.291790140808977e+17, 1.291790140849603e+17, 1.291790140890226e+17, 1.291790140932415e+17, 1.291790140971478e+17, 1.291790141012101e+17, 1.291790141052727e+17, 1.291790141093352e+17, 1.291790141133976e+17, 1.291790141174602e+17, 1.291790141215227e+17, 1.291790141255852e+17, 1.291790141296476e+17, 1.291790141337102e+17, 1.291790141377727e+17, 1.291790141418351e+17, 1.291790141458976e+17, 1.291790141499602e+17, 1.291790141540227e+17, 1.291790141580852e+17, 1.291790141621477e+17, 1.291790141662102e+17, 1.291790141702726e+17, 1.291790141743352e+17, 1.291790141783976e+17, 1.291790141824602e+17, 1.291790141865228e+17, 1.291790141905851e+17, 1.291790141946477e+17, 1.291790141987103e+17, 1.291790142027727e+17, 1.291790142068351e+17, 1.291790142108977e+17, 1.291790142149603e+17, 1.291790142190227e+17, 1.291790142230852e+17, 1.291790142271476e+17, 1.291790142312101e+17, 1.291790142352727e+17, 1.291790142393352e+17, 1.291790142433976e+17, 1.291790142476164e+17, 1.291790142515227e+17, 1.291790142555852e+17, 1.291790142596476e+17, 1.291790142637102e+17, 1.291790142677727e+17, 1.291790142718351e+17, 1.291790142760539e+17, 1.291790142799602e+17, 1.291790142840227e+17, 1.291790142880851e+17, 1.291790142921477e+17, 1.291790142962102e+17, 1.291790143002726e+17, 1.291790143043352e+17, 1.291790143083976e+17, 1.291790143124602e+17, 1.291790143165228e+17, 1.291790143205851e+17, 1.291790143246477e+17, 1.291790143287101e+17, 1.291790143327727e+17, 1.291790143368352e+17, 1.291790143408977e+17, 1.291790143449603e+17, 1.291790143490226e+17, 1.291790143530852e+17, 1.291790143571478e+17, 1.291790143612101e+17, 1.291790143652727e+17, 1.291790143693352e+17, 1.291790143735539e+17, 1.291790143774602e+17, 1.291790143815227e+17, 1.291790143855852e+17, 1.291790143896476e+17, 1.291790143937102e+17, 1.291790143977727e+17, 1.291790144018351e+17, 1.291790144058976e+17, 1.291790144099602e+17, 1.291790144140227e+17, 1.291790144180852e+17, 1.291790144221477e+17, 1.291790144262102e+17, 1.291790144302726e+17, 1.291790144343352e+17, 1.291790144383976e+17, 1.291790144424602e+17, 1.291790144465228e+17, 1.291790144505851e+17, 1.291790144546477e+17, 1.291790144587103e+17, 1.291790144627726e+17, 1.291790144668352e+17, 1.291790144708977e+17, 1.291790144749603e+17, 1.291790144790227e+17, 1.291790144830852e+17, 1.291790144871476e+17, 1.291790144912101e+17, 1.291790144952727e+17, 1.291790144993353e+17, 1.291790145033976e+17, 1.291790145074601e+17, 1.291790145115227e+17, 1.291790145155852e+17, 1.291790145196476e+17, 1.291790145237102e+17, 1.291790145277727e+17, 1.291790145316788e+17, 1.291790145358977e+17, 1.291790145399602e+17, 1.291790145440227e+17, 1.291790145480851e+17, 1.291790145519914e+17, 1.291790145562102e+17, 1.291790145602726e+17, 1.291790145643352e+17, 1.291790145683976e+17, 1.291790145724602e+17, 1.291790145765228e+17, 1.291790145805851e+17, 1.291790145846477e+17, 1.291790145887101e+17, 1.291790145927726e+17, 1.291790145968352e+17, 1.291790146008977e+17, 1.291790146049601e+17, 1.291790146090226e+17, 1.291790146130852e+17, 1.291790146171478e+17, 1.291790146212101e+17, 1.291790146252727e+17, 1.291790146293352e+17, 1.291790146333976e+17, 1.291790146374602e+17, 1.291790146415227e+17, 1.291790146455852e+17, 1.291790146496476e+17, 1.291790146537102e+17, 1.291790146577727e+17, 1.291790146618351e+17, 1.291790146658976e+17, 1.291790146699602e+17, 1.291790146740227e+17, 1.291790146780852e+17, 1.291790146821477e+17, 1.291790146862102e+17, 1.291790146902726e+17, 1.291790146943352e+17, 1.291790146983976e+17, 1.291790147024602e+17, 1.291790147065228e+17, 1.291790147105851e+17, 1.291790147146477e+17, 1.291790147187103e+17, 1.291790147227726e+17, 1.291790147268352e+17, 1.291790147308977e+17, 1.291790147349601e+17, 1.291790147390227e+17, 1.291790147430852e+17, 1.291790147471476e+17, 1.291790147512101e+17, 1.291790147552727e+17, 1.291790147591789e+17, 1.291790147633976e+17, 1.291790147674601e+17, 1.291790147715227e+17, 1.291790147755852e+17, 1.291790147796476e+17, 1.291790147837102e+17, 1.291790147877727e+17, 1.291790147918351e+17, 1.291790147958977e+17, 1.291790147999602e+17, 1.291790148040227e+17, 1.291790148080851e+17, 1.291790148121477e+17, 1.291790148162102e+17, 1.291790148202726e+17, 1.291790148243352e+17, 1.291790148283976e+17, 1.291790148324602e+17, 1.291790148365228e+17, 1.291790148405851e+17, 1.291790148446477e+17, 1.291790148487101e+17, 1.291790148527726e+17, 1.291790148568352e+17, 1.291790148608977e+17, 1.291790148649601e+17, 1.291790148690226e+17, 1.291790148730852e+17, 1.291790148771476e+17, 1.291790148812101e+17, 1.291790148852727e+17, 1.291790148893352e+17, 1.291790148933976e+17, 1.291790148974602e+17, 1.291790149015227e+17, 1.291790149055852e+17, 1.291790149096476e+17, 1.291790149137102e+17, 1.291790149177727e+17, 1.291790149218351e+17, 1.291790149258976e+17, 1.291790149299602e+17, 1.291790149340227e+17, 1.291790149380852e+17, 1.291790149421477e+17, 1.291790149462102e+17, 1.291790149502726e+17, 1.291790149543352e+17, 1.291790149583976e+17, 1.291790149624602e+17, 1.291790149665228e+17, 1.291790149705851e+17, 1.291790149746477e+17, 1.291790149787103e+17, 1.291790149827726e+17, 1.291790149868352e+17, 1.291790149908977e+17, 1.291790149949601e+17, 1.291790149990227e+17, 1.291790150030852e+17, 1.291790150071476e+17, 1.291790150112101e+17, 1.291790150152727e+17, 1.291790150193353e+17, 1.291790150233976e+17, 1.291790150274601e+17, 1.291790150315227e+17, 1.291790150355852e+17, 1.291790150396476e+17, 1.291790150437102e+17, 1.291790150477727e+17, 1.291790150518351e+17, 1.291790150558977e+17, 1.291790150599602e+17, 1.291790150640227e+17, 1.291790150680851e+17, 1.291790150721477e+17, 1.291790150762102e+17, 1.291790150802726e+17, 1.291790150843352e+17, 1.291790150883976e+17, 1.291790150924602e+17, 1.291790150965228e+17, 1.291790151005851e+17, 1.291790151046477e+17, 1.291790151087101e+17, 1.291790151127726e+17, 1.291790151168352e+17, 1.291790151208977e+17, 1.291790151249601e+17, 1.291790151290226e+17, 1.291790151330852e+17, 1.291790151371476e+17, 1.291790151412101e+17, 1.291790151452727e+17, 1.291790151493352e+17, 1.291790151533976e+17, 1.291790151574602e+17, 1.291790151615227e+17, 1.291790151655852e+17, 1.291790151696476e+17, 1.291790151737102e+17, 1.291790151777727e+17, 1.291790151818351e+17, 1.291790151858976e+17, 1.291790151899602e+17, 1.291790151940227e+17, 1.291790151980852e+17, 1.291790152021477e+17, 1.291790152062102e+17, 1.291790152102726e+17, 1.291790152143352e+17, 1.291790152183976e+17, 1.291790152224602e+17, 1.291790152265228e+17, 1.291790152305851e+17, 1.291790152346477e+17, 1.291790152387103e+17, 1.291790152427726e+17, 1.291790152468352e+17, 1.291790152508977e+17, 1.291790152549601e+17, 1.291790152590227e+17, 1.291790152630852e+17, 1.291790152671476e+17, 1.291790152712101e+17, 1.291790152752727e+17, 1.291790152793352e+17, 1.291790152833976e+17, 1.291790152874602e+17, 1.291790152915227e+17, 1.291790152955852e+17, 1.291790152996476e+17, 1.291790153037102e+17, 1.291790153077727e+17, 1.291790153118351e+17, 1.291790153158977e+17, 1.291790153199602e+17, 1.291790153240227e+17, 1.291790153280851e+17, 1.291790153321477e+17, 1.291790153362102e+17, 1.291790153402726e+17, 1.291790153444914e+17, 1.29179015348554e+17, 1.291790153524602e+17, 1.291790153565228e+17, 1.291790153605851e+17, 1.291790153646477e+17, 1.291790153687101e+17, 1.291790153727726e+17, 1.291790153768352e+17, 1.291790153808977e+17, 1.291790153849601e+17, 1.291790153890226e+17, 1.291790153930852e+17, 1.291790153971476e+17, 1.291790154012101e+17, 1.291790154052727e+17, 1.291790154093352e+17, 1.291790154133976e+17, 1.291790154174602e+17, 1.291790154215227e+17, 1.291790154255852e+17, 1.291790154296476e+17, 1.291790154337102e+17, 1.291790154377727e+17, 1.291790154418351e+17, 1.291790154458976e+17, 1.291790154499602e+17, 1.291790154540227e+17, 1.291790154580852e+17, 1.291790154621477e+17, 1.291790154662102e+17, 1.291790154702726e+17, 1.291790154743352e+17, 1.291790154783976e+17, 1.291790154824602e+17, 1.291790154865228e+17, 1.291790154905851e+17, 1.291790154946477e+17, 1.291790154987103e+17, 1.291790155027726e+17, 1.291790155068352e+17, 1.291790155108977e+17, 1.291790155149601e+17, 1.291790155190227e+17, 1.291790155230852e+17, 1.291790155271476e+17, 1.291790155312101e+17, 1.291790155352727e+17, 1.291790155393352e+17, 1.291790155433976e+17, 1.291790155474602e+17, 1.291790155515227e+17, 1.291790155555852e+17, 1.291790155596476e+17, 1.291790155637102e+17, 1.291790155677727e+17, 1.291790155718351e+17, 1.291790155758977e+17, 1.291790155799602e+17, 1.291790155840227e+17, 1.291790155880851e+17, 1.291790155921477e+17, 1.291790155962102e+17, 1.291790156002726e+17, 1.291790156043352e+17, 1.291790156083976e+17, 1.291790156124602e+17, 1.291790156165228e+17, 1.291790156205851e+17, 1.291790156246477e+17, 1.291790156287101e+17, 1.291790156327726e+17, 1.291790156368352e+17, 1.291790156408977e+17, 1.291790156449601e+17, 1.291790156490226e+17, 1.291790156530852e+17, 1.291790156571476e+17, 1.291790156612101e+17, 1.291790156652727e+17, 1.291790156691789e+17, 1.291790156733976e+17, 1.291790156774602e+17, 1.291790156815227e+17, 1.291790156855852e+17, 1.291790156896476e+17, 1.291790156937102e+17, 1.291790156977727e+17, 1.291790157018351e+17, 1.291790157058977e+17, 1.291790157099602e+17, 1.291790157140227e+17, 1.291790157180852e+17, 1.291790157221477e+17, 1.291790157262102e+17, 1.291790157302726e+17, 1.291790157343352e+17, 1.291790157383977e+17, 1.291790157424602e+17, 1.291790157465228e+17, 1.291790157505851e+17, 1.291790157546477e+17, 1.291790157587103e+17, 1.291790157627726e+17, 1.291790157668352e+17, 1.291790157708977e+17, 1.291790157749601e+17, 1.291790157790227e+17, 1.291790157830852e+17, 1.291790157871476e+17, 1.291790157912101e+17, 1.291790157952727e+17, 1.291790157993352e+17, 1.291790158033976e+17, 1.291790158074602e+17, 1.291790158115227e+17, 1.291790158155852e+17, 1.291790158196476e+17, 1.291790158237102e+17, 1.291790158277727e+17, 1.291790158318351e+17, 1.291790158358977e+17, 1.291790158399602e+17, 1.291790158440227e+17, 1.291790158480851e+17, 1.291790158521477e+17, 1.291790158562102e+17, 1.291790158602728e+17, 1.291790158643352e+17, 1.291790158683976e+17, 1.291790158724602e+17, 1.291790158765228e+17, 1.291790158805851e+17, 1.291790158846477e+17, 1.291790158887101e+17, 1.291790158927726e+17, 1.291790158969914e+17, 1.291790159008977e+17, 1.291790159049601e+17, 1.291790159090226e+17, 1.291790159130852e+17, 1.291790159171476e+17, 1.291790159212101e+17, 1.291790159252727e+17, 1.291790159293352e+17, 1.291790159333976e+17, 1.291790159374602e+17, 1.291790159415227e+17, 1.291790159455852e+17, 1.291790159496476e+17, 1.291790159537102e+17, 1.291790159577727e+17, 1.291790159618351e+17, 1.291790159658977e+17, 1.291790159699602e+17, 1.291790159740227e+17, 1.291790159780852e+17, 1.291790159821477e+17, 1.291790159862102e+17, 1.291790159902726e+17, 1.291790159943352e+17, 1.291790159983977e+17, 1.291790160024602e+17, 1.291790160065228e+17, 1.291790160105851e+17, 1.291790160146477e+17, 1.291790160187103e+17, 1.291790160227726e+17, 1.291790160268352e+17, 1.291790160308977e+17, 1.291790160349601e+17, 1.291790160390227e+17, 1.291790160430852e+17, 1.291790160471476e+17, 1.291790160513664e+17, 1.291790160554289e+17, 1.291790160594915e+17, 1.291790160633976e+17, 1.291790160676164e+17, 1.291790160715227e+17, 1.291790160755852e+17, 1.291790160796476e+17, 1.291790160837102e+17, 1.291790160877727e+17, 1.291790160918351e+17, 1.291790160958977e+17, 1.291790160999602e+17, 1.291790161040227e+17, 1.291790161080852e+17, 1.291790161121477e+17, 1.291790161162102e+17, 1.291790161202728e+17, 1.291790161243352e+17, 1.291790161283976e+17, 1.291790161324602e+17, 1.291790161365228e+17, 1.291790161405852e+17, 1.291790161446477e+17, 1.291790161487101e+17, 1.29179016152929e+17, 1.291790161569914e+17, 1.29179016161054e+17, 1.291790161651164e+17, 1.291790161690226e+17, 1.291790161730852e+17, 1.291790161771476e+17, 1.291790161812101e+17, 1.291790161852727e+17, 1.291790161893352e+17, 1.291790161933976e+17, 1.291790161974602e+17, 1.291790162015227e+17, 1.291790162055852e+17, 1.291790162096476e+17, 1.291790162137102e+17, 1.291790162177727e+17, 1.291790162218351e+17, 1.291790162258977e+17, 1.291790162299602e+17, 1.291790162340227e+17, 1.291790162380852e+17, 1.291790162421477e+17, 1.291790162462102e+17, 1.291790162502726e+17, 1.291790162543352e+17, 1.291790162583977e+17, 1.291790162624602e+17, 1.291790162665228e+17, 1.291790162705851e+17, 1.291790162746477e+17, 1.291790162787103e+17, 1.291790162827726e+17, 1.291790162868352e+17, 1.291790162908977e+17, 1.291790162949601e+17, 1.291790162990227e+17, 1.291790163030852e+17, 1.291790163071476e+17, 1.291790163112101e+17, 1.291790163152727e+17, 1.291790163193352e+17, 1.291790163233976e+17, 1.291790163274602e+17, 1.291790163315227e+17, 1.291790163355852e+17, 1.291790163396476e+17, 1.291790163437102e+17, 1.291790163477727e+17, 1.291790163518351e+17, 1.291790163558977e+17, 1.291790163599602e+17, 1.291790163640227e+17, 1.291790163680852e+17, 1.291790163721477e+17, 1.291790163762102e+17, 1.291790163802728e+17, 1.291790163843352e+17, 1.291790163883976e+17, 1.291790163924602e+17, 1.291790163965228e+17, 1.291790164005852e+17, 1.291790164046477e+17, 1.291790164087101e+17, 1.291790164127726e+17, 1.291790164168352e+17, 1.291790164208977e+17, 1.291790164249601e+17, 1.291790164290226e+17, 1.291790164330852e+17, 1.291790164371476e+17, 1.291790164412101e+17, 1.291790164452727e+17, 1.291790164493352e+17, 1.291790164533976e+17, 1.291790164574602e+17, 1.291790164615227e+17, 1.291790164655852e+17, 1.291790164696476e+17, 1.291790164737102e+17, 1.291790164777727e+17, 1.291790164818351e+17, 1.291790164858977e+17, 1.291790164899601e+17, 1.291790164940227e+17, 1.291790164980852e+17, 1.291790165019914e+17, 1.291790165062102e+17, 1.291790165102726e+17, 1.291790165143352e+17, 1.291790165183977e+17, 1.291790165224602e+17, 1.291790165265228e+17, 1.291790165305851e+17, 1.291790165346477e+17, 1.291790165387103e+17, 1.291790165427726e+17, 1.291790165468352e+17, 1.291790165508977e+17, 1.291790165549601e+17, 1.291790165590227e+17, 1.291790165630852e+17, 1.291790165671476e+17, 1.291790165712101e+17, 1.291790165752727e+17, 1.291790165793352e+17, 1.291790165833976e+17, 1.291790165874602e+17, 1.291790165915227e+17, 1.291790165955852e+17, 1.291790165996476e+17, 1.291790166037102e+17, 1.291790166077727e+17, 1.291790166118351e+17, 1.291790166158977e+17, 1.291790166199602e+17, 1.291790166240227e+17, 1.291790166280852e+17, 1.291790166321476e+17, 1.291790166362102e+17, 1.291790166402728e+17, 1.291790166443352e+17, 1.291790166483976e+17, 1.291790166524602e+17, 1.291790166565228e+17, 1.291790166605852e+17, 1.291790166646477e+17, 1.291790166687101e+17, 1.291790166727726e+17, 1.291790166768352e+17, 1.291790166808977e+17, 1.291790166849601e+17, 1.291790166890226e+17, 1.291790166929289e+17, 1.291790166971476e+17, 1.291790167012101e+17, 1.291790167052727e+17, 1.291790167093352e+17, 1.291790167133976e+17, 1.291790167174602e+17, 1.291790167215227e+17, 1.291790167255852e+17, 1.291790167296476e+17, 1.291790167337102e+17, 1.291790167377727e+17, 1.291790167418351e+17, 1.291790167458977e+17, 1.291790167499601e+17, 1.291790167540227e+17, 1.291790167580852e+17, 1.291790167621476e+17, 1.291790167662102e+17, 1.291790167702726e+17, 1.291790167743352e+17, 1.291790167783977e+17, 1.291790167824602e+17, 1.291790167865228e+17, 1.291790167905851e+17, 1.29179016794804e+17, 1.291790167988664e+17, 1.291790168027726e+17, 1.291790168068352e+17, 1.291790168108977e+17, 1.291790168149601e+17, 1.291790168190227e+17, 1.291790168230852e+17, 1.291790168271476e+17, 1.291790168312101e+17, 1.291790168352727e+17, 1.291790168393352e+17, 1.291790168433976e+17, 1.291790168474602e+17, 1.291790168515227e+17, 1.291790168555852e+17, 1.291790168596476e+17, 1.291790168637102e+17, 1.291790168677727e+17, 1.291790168718351e+17, 1.291790168758977e+17, 1.291790168799602e+17, 1.291790168840227e+17, 1.291790168880852e+17, 1.291790168921476e+17, 1.291790168962102e+17, 1.291790169002728e+17, 1.291790169043351e+17, 1.291790169083976e+17, 1.291790169124602e+17, 1.291790169165228e+17, 1.291790169205852e+17, 1.291790169246477e+17, 1.291790169287103e+17, 1.291790169327726e+17, 1.291790169368352e+17, 1.291790169408977e+17, 1.29179016944804e+17, 1.291790169490226e+17, 1.291790169530852e+17, 1.291790169571476e+17, 1.291790169612102e+17, 1.291790169652727e+17, 1.291790169693352e+17, 1.291790169733976e+17, 1.291790169774602e+17, 1.291790169815227e+17, 1.291790169855852e+17, 1.291790169896476e+17, 1.291790169937102e+17, 1.291790169977727e+17, 1.29179017001679e+17, 1.291790170058977e+17, 1.291790170099601e+17, 1.291790170140227e+17, 1.291790170180852e+17, 1.291790170221476e+17, 1.291790170262102e+17, 1.291790170302726e+17, 1.291790170341788e+17, 1.291790170383977e+17, 1.291790170424602e+17, 1.291790170465228e+17, 1.291790170505851e+17, 1.291790170546477e+17, 1.291790170585539e+17, 1.291790170627726e+17, 1.291790170668352e+17, 1.291790170708977e+17, 1.291790170749601e+17, 1.291790170790227e+17, 1.291790170830852e+17, 1.291790170871476e+17, 1.291790170912101e+17, 1.291790170952727e+17, 1.291790170993352e+17, 1.291790171033976e+17, 1.291790171074602e+17, 1.291790171115227e+17, 1.291790171155852e+17, 1.291790171198039e+17, 1.291790171237102e+17, 1.291790171277727e+17, 1.291790171318351e+17, 1.291790171358977e+17, 1.291790171399602e+17, 1.291790171440227e+17, 1.29179017147929e+17, 1.291790171521476e+17, 1.291790171562102e+17, 1.291790171602728e+17, 1.291790171643351e+17, 1.291790171683976e+17, 1.291790171724602e+17, 1.291790171765226e+17, 1.291790171805852e+17, 1.291790171846477e+17, 1.291790171887103e+17, 1.291790171927726e+17, 1.291790171968352e+17, 1.291790172008977e+17, 1.291790172049601e+17, 1.291790172090227e+17, 1.291790172130852e+17, 1.291790172173039e+17, 1.291790172212102e+17, 1.291790172252727e+17, 1.291790172293352e+17, 1.291790172333976e+17, 1.291790172374602e+17, 1.291790172415227e+17, 1.291790172455852e+17, 1.291790172496476e+17, 1.291790172537102e+17, 1.291790172577727e+17, 1.291790172618351e+17, 1.291790172658977e+17, 1.291790172699601e+17, 1.291790172740227e+17, 1.291790172780852e+17, 1.291790172821476e+17, 1.291790172862102e+17, 1.291790172902726e+17, 1.291790172943351e+17, 1.291790172983977e+17, 1.291790173024602e+17, 1.291790173065226e+17, 1.291790173105851e+17, 1.291790173146477e+17, 1.291790173187101e+17, 1.291790173227726e+17, 1.291790173268352e+17, 1.291790173308977e+17, 1.291790173349601e+17, 1.291790173390227e+17, 1.291790173429289e+17, 1.291790173471476e+17, 1.291790173512101e+17, 1.291790173552727e+17, 1.291790173593352e+17, 1.291790173633976e+17, 1.291790173674602e+17, 1.291790173715227e+17, 1.291790173755852e+17, 1.291790173796477e+17, 1.291790173837102e+17, 1.291790173877727e+17, 1.291790173918351e+17, 1.291790173958977e+17, 1.291790173999602e+17, 1.291790174040227e+17, 1.291790174080852e+17, 1.291790174121476e+17, 1.291790174162102e+17, 1.291790174202728e+17, 1.291790174243351e+17, 1.291790174283976e+17, 1.291790174324602e+17, 1.291790174365226e+17, 1.291790174405852e+17, 1.291790174446477e+17, 1.291790174487101e+17, 1.291790174527726e+17, 1.291790174568352e+17, 1.291790174608977e+17, 1.291790174649601e+17, 1.291790174690227e+17, 1.291790174730852e+17, 1.291790174771476e+17, 1.291790174812102e+17, 1.291790174852727e+17, 1.291790174893352e+17, 1.291790174933976e+17, 1.291790174974602e+17, 1.291790175015227e+17, 1.291790175055852e+17, 1.291790175096476e+17, 1.291790175137102e+17, 1.291790175177727e+17, 1.291790175218351e+17, 1.291790175258977e+17, 1.291790175299601e+17, 1.291790175340227e+17, 1.291790175380852e+17, 1.291790175421476e+17, 1.291790175462102e+17, 1.291790175502726e+17, 1.291790175543351e+17, 1.291790175583977e+17, 1.291790175624602e+17, 1.291790175665226e+17, 1.291790175705851e+17, 1.291790175746477e+17, 1.291790175787101e+17, 1.291790175827726e+17, 1.291790175868352e+17, 1.291790175908977e+17, 1.291790175949601e+17, 1.291790175990227e+17, 1.291790176029289e+17, 1.291790176071476e+17, 1.291790176112101e+17, 1.291790176152727e+17, 1.291790176193352e+17, 1.291790176233976e+17, 1.291790176274602e+17, 1.291790176315227e+17, 1.291790176355852e+17, 1.291790176396477e+17, 1.291790176437102e+17, 1.291790176477727e+17, 1.291790176518351e+17, 1.291790176558977e+17, 1.291790176599602e+17, 1.291790176640227e+17, 1.291790176680852e+17, 1.291790176721476e+17, 1.291790176762102e+17, 1.291790176802728e+17, 1.291790176841789e+17, 1.291790176883976e+17, 1.291790176924602e+17, 1.291790176965226e+17, 1.291790177005852e+17, 1.291790177046477e+17, 1.291790177087101e+17, 1.291790177127726e+17, 1.291790177168352e+17, 1.291790177208977e+17, 1.291790177249601e+17, 1.291790177290227e+17, 1.291790177330852e+17, 1.291790177371476e+17, 1.291790177412102e+17, 1.291790177452727e+17, 1.291790177493352e+17, 1.291790177533976e+17, 1.291790177574602e+17, 1.291790177615227e+17, 1.291790177655852e+17, 1.291790177696476e+17, 1.291790177737102e+17, 1.291790177777727e+17, 1.291790177818353e+17, 1.291790177858977e+17, 1.291790177899601e+17, 1.291790177940227e+17, 1.291790177980852e+17, 1.291790178021476e+17, 1.291790178062102e+17, 1.291790178102726e+17, 1.291790178143351e+17, 1.291790178183977e+17, 1.291790178224602e+17, 1.291790178265226e+17, 1.291790178305851e+17, 1.291790178346477e+17, 1.291790178387101e+17, 1.291790178427726e+17, 1.291790178468352e+17, 1.291790178508977e+17, 1.291790178549601e+17, 1.291790178590227e+17, 1.291790178630852e+17, 1.291790178671476e+17, 1.291790178712101e+17, 1.291790178752727e+17, 1.291790178793352e+17, 1.291790178833976e+17, 1.291790178874602e+17, 1.291790178915227e+17, 1.291790178955852e+17, 1.291790178996477e+17, 1.291790179037102e+17, 1.291790179077727e+17, 1.291790179118351e+17, 1.291790179158977e+17, 1.291790179199602e+17, 1.291790179240227e+17, 1.291790179280852e+17, 1.291790179321476e+17, 1.291790179362102e+17, 1.291790179402728e+17, 1.291790179443351e+17, 1.291790179483976e+17, 1.291790179524602e+17, 1.291790179565226e+17, 1.291790179605852e+17, 1.291790179646477e+17, 1.291790179685539e+17, 1.291790179727726e+17, 1.291790179768352e+17, 1.291790179808977e+17, 1.291790179849601e+17, 1.291790179890227e+17, 1.291790179930852e+17, 1.291790179971476e+17, 1.291790180012102e+17, 1.291790180052727e+17, 1.291790180093352e+17, 1.291790180133976e+17, 1.291790180174602e+17, 1.291790180215227e+17, 1.29179018025429e+17, 1.291790180296476e+17, 1.291790180337102e+17, 1.291790180377727e+17, 1.291790180418353e+17, 1.291790180458977e+17, 1.291790180499601e+17, 1.291790180540227e+17, 1.291790180579288e+17, 1.291790180621476e+17, 1.291790180662102e+17, 1.291790180702726e+17, 1.291790180743351e+17, 1.291790180783977e+17, 1.291790180824602e+17, 1.291790180865226e+17, 1.291790180905851e+17, 1.291790180946477e+17, 1.291790180987101e+17, 1.291790181027726e+17, 1.291790181068352e+17, 1.291790181108977e+17, 1.291790181149601e+17, 1.291790181190227e+17, 1.291790181230852e+17, 1.291790181271476e+17, 1.291790181312101e+17, 1.291790181352727e+17, 1.291790181393352e+17, 1.291790181433976e+17, 1.291790181474602e+17, 1.291790181515227e+17, 1.291790181555852e+17, 1.291790181596477e+17, 1.291790181637102e+17, 1.291790181677727e+17, 1.29179018171679e+17, 1.291790181758977e+17, 1.291790181799602e+17, 1.291790181840227e+17, 1.291790181880852e+17, 1.291790181921476e+17, 1.291790181962102e+17, 1.291790182002728e+17, 1.291790182043351e+17, 1.291790182083976e+17, 1.291790182124602e+17, 1.291790182165226e+17, 1.291790182205852e+17, 1.291790182246477e+17, 1.291790182287101e+17, 1.291790182327726e+17, 1.291790182368352e+17, 1.291790182408977e+17, 1.291790182449601e+17, 1.291790182490227e+17, 1.291790182530852e+17, 1.291790182571476e+17, 1.291790182612102e+17, 1.291790182652727e+17, 1.291790182693352e+17, 1.291790182733976e+17, 1.291790182774602e+17, 1.291790182815227e+17, 1.291790182855852e+17, 1.291790182896476e+17, 1.291790182937102e+17, 1.291790182977727e+17, 1.291790183018353e+17, 1.291790183058977e+17, 1.291790183099601e+17, 1.291790183140227e+17, 1.291790183180852e+17, 1.291790183221476e+17, 1.291790183262102e+17, 1.291790183302726e+17, 1.291790183343351e+17, 1.291790183383977e+17, 1.291790183424602e+17, 1.291790183465226e+17, 1.291790183505851e+17, 1.291790183546477e+17, 1.291790183587101e+17, 1.291790183627726e+17, 1.291790183668352e+17, 1.291790183708977e+17, 1.291790183749601e+17, 1.291790183790227e+17, 1.291790183830852e+17, 1.291790183871476e+17, 1.291790183912101e+17, 1.291790183952727e+17, 1.291790183993352e+17, 1.291790184033976e+17, 1.291790184074602e+17, 1.291790184115227e+17, 1.291790184155852e+17, 1.291790184196477e+17, 1.291790184237102e+17, 1.291790184277727e+17, 1.291790184318351e+17, 1.291790184358977e+17, 1.291790184399602e+17, 1.291790184440227e+17, 1.291790184480852e+17, 1.291790184521476e+17, 1.291790184562102e+17, 1.291790184602728e+17, 1.291790184643351e+17, 1.291790184683976e+17, 1.291790184724602e+17, 1.291790184765226e+17, 1.291790184804289e+17, 1.291790184844914e+17, 1.291790184887101e+17, 1.291790184927726e+17, 1.291790184968352e+17, 1.291790185008977e+17, 1.291790185049601e+17, 1.291790185090227e+17, 1.291790185130852e+17, 1.291790185171476e+17, 1.291790185212102e+17, 1.291790185252727e+17, 1.291790185293352e+17, 1.291790185333976e+17, 1.291790185374602e+17, 1.291790185415227e+17, 1.291790185455852e+17, 1.291790185496476e+17, 1.291790185537102e+17, 1.291790185577727e+17, 1.291790185618353e+17, 1.291790185658977e+17, 1.291790185699602e+17, 1.291790185740227e+17, 1.291790185780852e+17, 1.291790185821476e+17, 1.291790185862102e+17, 1.291790185902726e+17, 1.291790185943351e+17, 1.291790185983977e+17, 1.291790186024603e+17, 1.291790186065226e+17, 1.291790186105851e+17, 1.291790186146477e+17, 1.291790186187101e+17, 1.291790186227726e+17, 1.291790186268352e+17, 1.291790186308977e+17, 1.291790186349601e+17, 1.291790186390227e+17, 1.291790186430852e+17, 1.291790186471476e+17, 1.291790186512101e+17, 1.291790186552727e+17, 1.291790186593352e+17, 1.291790186633976e+17, 1.291790186674602e+17, 1.291790186715227e+17, 1.291790186755852e+17, 1.291790186796477e+17, 1.291790186837102e+17, 1.291790186877727e+17, 1.291790186918351e+17, 1.291790186958977e+17, 1.291790186999602e+17, 1.291790187040227e+17, 1.291790187080852e+17, 1.291790187121476e+17, 1.291790187162102e+17, 1.291790187202728e+17, 1.291790187243351e+17, 1.291790187283976e+17, 1.291790187324602e+17, 1.291790187365226e+17, 1.291790187405852e+17, 1.291790187446477e+17, 1.291790187487101e+17, 1.291790187527726e+17, 1.291790187568352e+17, 1.291790187608977e+17, 1.291790187649601e+17, 1.291790187690227e+17, 1.291790187730852e+17, 1.291790187771476e+17, 1.291790187812102e+17, 1.291790187852727e+17, 1.291790187893352e+17, 1.291790187933976e+17, 1.291790187974602e+17, 1.291790188015227e+17, 1.291790188055852e+17, 1.291790188096476e+17, 1.291790188137102e+17, 1.291790188177727e+17, 1.291790188218353e+17, 1.291790188258977e+17, 1.291790188299602e+17, 1.291790188340227e+17, 1.291790188380852e+17, 1.291790188421476e+17, 1.291790188462102e+17, 1.291790188502728e+17, 1.291790188543351e+17, 1.291790188583977e+17, 1.291790188624603e+17, 1.291790188665226e+17, 1.291790188705851e+17, 1.291790188746477e+17, 1.291790188785539e+17, 1.291790188827727e+17, 1.291790188868352e+17, 1.291790188908977e+17, 1.291790188949601e+17, 1.291790188990227e+17, 1.291790189030852e+17, 1.291790189071476e+17, 1.291790189112101e+17, 1.291790189152727e+17, 1.291790189193352e+17, 1.291790189233976e+17, 1.291790189274602e+17, 1.291790189315226e+17, 1.291790189355852e+17, 1.291790189396477e+17, 1.291790189437102e+17, 1.291790189477727e+17, 1.291790189518351e+17, 1.291790189558977e+17, 1.291790189599602e+17, 1.291790189640227e+17, 1.29179018967929e+17, 1.291790189721476e+17, 1.291790189762102e+17, 1.291790189802728e+17, 1.291790189843351e+17, 1.291790189883977e+17, 1.291790189924602e+17, 1.291790189966789e+17, 1.291790190005852e+17, 1.291790190046477e+17, 1.291790190087101e+17, 1.291790190127726e+17, 1.291790190168352e+17, 1.291790190208977e+17, 1.291790190249601e+17, 1.291790190290227e+17, 1.291790190330852e+17, 1.291790190371476e+17, 1.291790190412102e+17, 1.291790190452727e+17, 1.291790190493352e+17, 1.291790190533976e+17, 1.291790190574602e+17, 1.291790190615227e+17, 1.291790190655852e+17, 1.291790190696476e+17, 1.291790190737101e+17, 1.291790190777727e+17, 1.291790190818353e+17, 1.291790190858977e+17, 1.291790190899602e+17, 1.291790190940227e+17, 1.291790190980852e+17, 1.291790191021476e+17, 1.291790191062102e+17, 1.291790191102728e+17, 1.291790191143351e+17, 1.291790191183977e+17, 1.291790191224603e+17, 1.291790191265226e+17, 1.291790191305852e+17, 1.291790191346477e+17, 1.291790191387101e+17, 1.291790191427727e+17, 1.291790191468352e+17, 1.291790191508977e+17, 1.291790191549601e+17, 1.291790191590227e+17, 1.291790191629289e+17, 1.291790191671476e+17, 1.291790191712101e+17, 1.291790191752727e+17, 1.291790191793352e+17, 1.291790191833976e+17, 1.291790191874602e+17, 1.291790191915226e+17, 1.291790191955852e+17, 1.291790191996477e+17, 1.291790192037101e+17, 1.291790192077727e+17, 1.291790192118351e+17, 1.291790192158977e+17, 1.291790192199602e+17, 1.291790192240227e+17, 1.291790192280852e+17, 1.291790192319914e+17, 1.291790192362102e+17, 1.291790192402728e+17, 1.291790192443351e+17, 1.291790192483977e+17, 1.291790192524602e+17, 1.291790192565226e+17, 1.291790192605852e+17, 1.291790192646477e+17, 1.291790192687101e+17, 1.291790192727726e+17, 1.291790192768352e+17, 1.291790192808977e+17, 1.291790192849601e+17, 1.291790192890227e+17, 1.291790192930852e+17, 1.291790192971476e+17, 1.291790193012102e+17, 1.291790193052727e+17, 1.291790193091789e+17, 1.291790193133976e+17, 1.291790193174602e+17, 1.291790193215227e+17, 1.291790193255852e+17, 1.291790193296476e+17, 1.291790193337101e+17, 1.291790193377727e+17, 1.291790193418353e+17, 1.291790193458976e+17, 1.291790193499602e+17, 1.291790193540227e+17, 1.291790193580852e+17, 1.291790193621476e+17, 1.291790193662102e+17, 1.291790193702728e+17, 1.291790193743351e+17, 1.291790193783977e+17, 1.291790193824603e+17, 1.291790193865226e+17, 1.291790193905852e+17, 1.291790193944914e+17, 1.291790193987101e+17, 1.291790194027727e+17, 1.291790194068352e+17, 1.291790194108977e+17, 1.291790194149601e+17, 1.291790194190227e+17, 1.291790194229289e+17, 1.291790194271476e+17, 1.291790194312101e+17, 1.291790194352727e+17, 1.291790194393352e+17, 1.291790194433976e+17, 1.291790194474602e+17, 1.291790194515226e+17, 1.291790194555852e+17, 1.291790194596477e+17, 1.291790194637101e+17, 1.291790194677727e+17, 1.291790194718351e+17, 1.291790194758976e+17, 1.291790194799602e+17, 1.291790194840227e+17, 1.291790194880852e+17, 1.291790194921476e+17, 1.291790194962102e+17, 1.291790195002728e+17, 1.291790195043351e+17, 1.291790195083977e+17, 1.291790195124602e+17, 1.291790195165226e+17, 1.291790195205852e+17, 1.291790195246477e+17, 1.291790195287101e+17, 1.291790195327726e+17, 1.291790195369915e+17},
			             {1.291790126387101e+17, 1.291790126427727e+17, 1.291790126468351e+17, 1.291790126508977e+17, 1.291790126549603e+17, 1.291790126590226e+17, 1.291790126630852e+17, 1.291790126671476e+17, 1.291790126712101e+17, 1.291790126752727e+17, 1.291790126793352e+17, 1.291790126833976e+17, 1.291790126874601e+17},
			             {1.291790101932415e+17, 1.291790101971476e+17, 1.291790102012102e+17, 1.291790102052726e+17, 1.291790102093352e+17, 1.291790102133978e+17, 1.291790102174601e+17, 1.291790102215227e+17, 1.291790102255852e+17, 1.291790102296476e+17, 1.291790102337102e+17, 1.291790102377727e+17, 1.291790102418351e+17, 1.291790102458976e+17, 1.291790102499602e+17, 1.291790102540227e+17, 1.291790102580851e+17, 1.291790102621476e+17, 1.291790102662102e+17, 1.291790102702726e+17, 1.291790102743352e+17, 1.291790102783977e+17},
			             {1.291790083244914e+17, 1.291790083283977e+17, 1.291790083324602e+17, 1.291790083365226e+17, 1.291790083405852e+17, 1.291790083446477e+17, 1.291790083487101e+17, 1.291790083527727e+17},
			             {1.291790109690227e+17, 1.291790109729289e+17, 1.291790109769915e+17, 1.291790109812102e+17, 1.291790109852726e+17, 1.291790109893352e+17, 1.291790109933978e+17, 1.291790109974601e+17},
			             {1.291790142840227e+17, 1.291790142880851e+17, 1.291790142921477e+17, 1.291790142962102e+17, 1.291790143002726e+17, 1.291790143043352e+17, 1.291790143083976e+17, 1.291790143124602e+17, 1.291790143165228e+17, 1.291790143205851e+17, 1.291790143246477e+17, 1.291790143287101e+17},
			             {1.291790136624602e+17, 1.291790136665226e+17, 1.291790136705852e+17, 1.291790136746477e+17, 1.291790136787103e+17, 1.291790136827727e+17, 1.291790136868351e+17, 1.291790136908977e+17, 1.291790136949603e+17, 1.291790136990226e+17},
			             {1.291790144505851e+17, 1.291790144546477e+17, 1.291790144587103e+17, 1.291790144627726e+17, 1.291790144668352e+17, 1.291790144708977e+17, 1.291790144749603e+17, 1.291790144790227e+17, 1.291790144830852e+17},
			             {1.291790122974602e+17, 1.291790123015227e+17, 1.291790123055852e+17, 1.291790123096476e+17, 1.291790123137102e+17, 1.291790123177727e+17, 1.291790123218351e+17, 1.291790123258976e+17},
			             {1.291790156368352e+17, 1.291790156408977e+17, 1.291790156449601e+17, 1.291790156490226e+17, 1.291790156530852e+17, 1.291790156571476e+17, 1.291790156612101e+17},
			             {1.291790190493352e+17, 1.291790190533976e+17, 1.291790190574602e+17, 1.291790190615227e+17, 1.291790190655852e+17, 1.291790190696476e+17, 1.291790190737101e+17, 1.291790190777727e+17, 1.291790190818353e+17, 1.291790190858977e+17, 1.291790190899602e+17, 1.291790190940227e+17, 1.291790190980852e+17, 1.291790191021476e+17, 1.291790191062102e+17, 1.291790191102728e+17, 1.291790191143351e+17, 1.291790191183977e+17, 1.291790191224603e+17, 1.291790191265226e+17, 1.291790191305852e+17},
			             {1.291790192077727e+17, 1.291790192118351e+17, 1.291790192158977e+17, 1.291790192199602e+17, 1.291790192240227e+17, 1.291790192280852e+17, 1.291790192319914e+17, 1.291790192362102e+17, 1.291790192402728e+17, 1.291790192443351e+17, 1.291790192483977e+17, 1.291790192524602e+17, 1.291790192565226e+17, 1.291790192605852e+17, 1.291790192646477e+17},
			             {1.291790192524602e+17, 1.291790192565226e+17, 1.291790192605852e+17, 1.291790192646477e+17, 1.291790192687101e+17, 1.291790192727726e+17, 1.291790192768352e+17, 1.291790192808977e+17, 1.291790192849601e+17, 1.291790192890227e+17, 1.291790192930852e+17, 1.291790192971476e+17, 1.291790193012102e+17, 1.291790193052727e+17, 1.291790193091789e+17, 1.291790193133976e+17, 1.291790193174602e+17, 1.291790193215227e+17, 1.291790193255852e+17, 1.291790193296476e+17, 1.291790193337101e+17, 1.291790193377727e+17, 1.291790193418353e+17, 1.291790193458976e+17, 1.291790193499602e+17, 1.291790193540227e+17, 1.291790193580852e+17, 1.291790193621476e+17, 1.291790193662102e+17, 1.291790193702728e+17, 1.291790193743351e+17, 1.291790193783977e+17, 1.291790193824603e+17, 1.291790193865226e+17, 1.291790193905852e+17, 1.291790193944914e+17, 1.291790193987101e+17, 1.291790194027727e+17, 1.291790194068352e+17, 1.291790194108977e+17, 1.291790194149601e+17, 1.291790194190227e+17, 1.291790194229289e+17, 1.291790194271476e+17, 1.291790194312101e+17},
			             {1.291790079180851e+17, 1.291790079221476e+17, 1.291790079262102e+17, 1.291790079302726e+17, 1.291790079343351e+17, 1.291790079383977e+17, 1.291790079424602e+17, 1.291790079465226e+17, 1.291790079505852e+17, 1.291790079546477e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
