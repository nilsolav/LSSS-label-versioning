netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 5;
			channels = 1;
			categories = 6;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0,  15.0, 248.1,  11.6,  51.1;
			max_depth =  451.5, 248.1, 456.3,  28.8, 225.0;
			start_time = 131315631974075776, 131315637639232000, 131315637639232000, 131315641114700672, 131315637650013184;
			end_time = 131315637639232000, 131315653102825728, 131315653102825728, 131315641145794432, 131315652261575808;
			region_id = 1, 2, 3, 4, 5;
			region_name = "Layer1","Layer2","Layer3","Layer1","Layer2";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "";
			region_category_names = "1", "6", "1", "6", "1", "6";
			region_category_proportions = 0.3, 0.7, 0.5, 0.5, 0.9, 0.1;
			region_category_ids = 1, 2, 3, 4, 5, 6;
			region_type = analysis, analysis, analysis, analysis, analysis;
			channel_names = "38";
			region_channels = 1, 1, 1;
			mask_times = {1.313156319740758e+17, 1.313156319851694e+17, 1.313156319953257e+17, 1.313156320056383e+17, 1.313156320162632e+17, 1.31315632026732e+17, 1.313156320370445e+17, 1.313156320476695e+17, 1.313156320587633e+17, 1.313156320689196e+17, 1.31315632079232e+17, 1.313156320897007e+17, 1.313156321000132e+17, 1.31315632110482e+17, 1.313156321211069e+17, 1.313156321314195e+17, 1.313156321415758e+17, 1.31315632152357e+17, 1.31315632162982e+17, 1.313156321736069e+17, 1.313156321837632e+17, 1.313156321940758e+17, 1.313156322045444e+17, 1.313156322151695e+17, 1.313156322256383e+17, 1.31315632236107e+17, 1.313156322472008e+17, 1.313156322573571e+17, 1.313156322673571e+17, 1.313156322781382e+17, 1.313156322889196e+17, 1.31315632299857e+17, 1.313156323100133e+17, 1.313156323201696e+17, 1.313156323306383e+17, 1.313156323412632e+17, 1.313156323517321e+17, 1.313156323625132e+17, 1.313156323728257e+17, 1.31315632382982e+17, 1.313156323931383e+17, 1.313156324031382e+17, 1.313156324136069e+17, 1.313156324240758e+17, 1.313156324351695e+17, 1.313156324453258e+17, 1.313156324564196e+17, 1.313156324670445e+17, 1.31315632479232e+17, 1.313156324895444e+17, 1.313156325007945e+17, 1.313156325109508e+17, 1.313156325214195e+17, 1.313156325320444e+17, 1.31315632542982e+17, 1.313156325531382e+17, 1.313156325634508e+17, 1.313156325740758e+17, 1.313156325843882e+17, 1.313156325951695e+17, 1.31315632605482e+17, 1.31315632616107e+17, 1.313156326268883e+17, 1.313156326373571e+17, 1.313156326481382e+17, 1.313156326597007e+17, 1.313156326701696e+17, 1.31315632680482e+17, 1.313156326912632e+17, 1.313156327020444e+17, 1.31315632712357e+17, 1.313156327226694e+17, 1.313156327331382e+17, 1.313156327439195e+17, 1.313156327539195e+17, 1.313156327645445e+17, 1.31315632774857e+17, 1.313156327853257e+17, 1.31315632796107e+17, 1.313156328062633e+17, 1.31315632816732e+17, 1.313156328276695e+17, 1.313156328384508e+17, 1.313156328487633e+17, 1.313156328589194e+17, 1.31315632869232e+17, 1.313156328795444e+17, 1.313156328897007e+17, 1.31315632900482e+17, 1.313156329114195e+17, 1.313156329217321e+17, 1.313156329326696e+17, 1.313156329434508e+17, 1.313156329540756e+17, 1.313156329643882e+17, 1.31315632974857e+17, 1.313156329862633e+17, 1.313156329976695e+17, 1.313156330076695e+17, 1.313156330176695e+17, 1.31315633028607e+17, 1.313156330389196e+17, 1.313156330495444e+17, 1.31315633059857e+17, 1.313156330701695e+17, 1.313156330807945e+17, 1.313156330912632e+17, 1.31315633101732e+17, 1.313156331123571e+17, 1.313156331234508e+17, 1.31315633133607e+17, 1.313156331440758e+17, 1.313156331542321e+17, 1.313156331651695e+17, 1.313156331762633e+17, 1.313156331865757e+17, 1.313156331968883e+17, 1.313156332073569e+17, 1.313156332176695e+17, 1.313156332278258e+17, 1.313156332384507e+17, 1.313156332489194e+17, 1.313156332595444e+17, 1.313156332701695e+17, 1.313156332803258e+17, 1.313156333003258e+17, 1.313156333115758e+17, 1.313156333225133e+17, 1.313156333340758e+17, 1.313156333450132e+17, 1.313156333557944e+17, 1.313156333673569e+17, 1.313156333779821e+17, 1.313156333979821e+17, 1.313156334082945e+17, 1.313156334184507e+17, 1.313156334384507e+17, 1.31315633449232e+17, 1.31315633460482e+17, 1.313156334707945e+17, 1.313156334809507e+17, 1.313156334911069e+17, 1.313156335012632e+17, 1.313156335118883e+17, 1.313156335222007e+17, 1.313156335322008e+17, 1.313156335426696e+17, 1.31315633553607e+17, 1.313156335640758e+17, 1.313156335742321e+17, 1.31315633584857e+17, 1.313156335953258e+17, 1.31315633605482e+17, 1.313156336156383e+17, 1.313156336262633e+17, 1.313156336368883e+17, 1.313156336472008e+17, 1.313156336575132e+17, 1.313156336678258e+17, 1.313156336782944e+17, 1.313156336889196e+17, 1.313156337001695e+17, 1.313156337103258e+17, 1.313156337203258e+17, 1.313156337314195e+17, 1.313156337422007e+17, 1.313156337528257e+17, 1.31315633763607e+17, 1.313156337740758e+17, 1.313156337851695e+17, 1.313156337957946e+17, 1.313156338062633e+17, 1.313156338165757e+17, 1.313156338276695e+17, 1.313156338378258e+17, 1.31315633847982e+17, 1.31315633858607e+17, 1.313156338690757e+17, 1.313156338797007e+17, 1.313156338900133e+17, 1.313156339007945e+17, 1.313156339112632e+17, 1.313156339214195e+17, 1.313156339315757e+17, 1.31315633941732e+17, 1.313156339522007e+17, 1.313156339625133e+17, 1.31315633972982e+17, 1.313156339832945e+17, 1.313156339937632e+17, 1.313156340042321e+17, 1.313156340147008e+17, 1.313156340256383e+17, 1.313156340359507e+17, 1.313156340459507e+17, 1.313156340562632e+17, 1.313156340668883e+17, 1.31315634077982e+17, 1.313156340881382e+17, 1.31315634099232e+17, 1.31315634109857e+17, 1.313156341203258e+17, 1.313156341315757e+17, 1.313156341415758e+17, 1.313156341520444e+17, 1.31315634162357e+17, 1.313156341728257e+17, 1.313156341832945e+17, 1.313156341940758e+17, 1.313156342047008e+17, 1.313156342147007e+17, 1.313156342256383e+17, 1.313156342362633e+17, 1.313156342470445e+17, 1.31315634257982e+17, 1.313156342681382e+17, 1.313156342782945e+17, 1.313156342889194e+17, 1.31315634299232e+17, 1.313156343101695e+17, 1.313156343209508e+17, 1.313156343312632e+17, 1.313156343415757e+17, 1.313156343525133e+17, 1.313156343631383e+17, 1.313156343737632e+17, 1.313156343839195e+17, 1.313156343939195e+17, 1.313156344042319e+17, 1.313156344150132e+17, 1.313156344250132e+17, 1.313156344353257e+17, 1.31315634445482e+17, 1.313156344564195e+17, 1.31315634466732e+17, 1.313156344768883e+17, 1.313156344879821e+17, 1.313156344981384e+17, 1.313156345082945e+17, 1.313156345193883e+17, 1.313156345297009e+17, 1.31315634539857e+17, 1.313156345501695e+17, 1.313156345603258e+17, 1.313156345718883e+17, 1.313156345825133e+17, 1.31315634592982e+17, 1.313156346031383e+17, 1.313156346137633e+17, 1.313156346240758e+17, 1.313156346347008e+17, 1.313156346453257e+17, 1.313156346556383e+17, 1.313156346665757e+17, 1.313156346778258e+17, 1.313156346881382e+17, 1.313156346989196e+17, 1.313156347090757e+17, 1.31315634719857e+17, 1.313156347300132e+17, 1.313156347403258e+17, 1.313156347515757e+17, 1.31315634762982e+17, 1.313156347737632e+17, 1.313156347843882e+17, 1.313156347945445e+17, 1.313156348059507e+17, 1.313156348162632e+17, 1.31315634826732e+17, 1.313156348368882e+17, 1.313156348476695e+17, 1.313156348578258e+17, 1.313156348678257e+17, 1.313156348787633e+17, 1.313156348895444e+17, 1.313156349001695e+17, 1.313156349103258e+17, 1.313156349209508e+17, 1.313156349318883e+17, 1.31315634942357e+17, 1.313156349528257e+17, 1.313156349631382e+17, 1.313156349742319e+17, 1.313156349845445e+17, 1.313156349951695e+17, 1.313156350053258e+17, 1.313156350159507e+17, 1.31315635026732e+17, 1.313156350378258e+17, 1.313156350479821e+17, 1.313156350582945e+17, 1.313156350684508e+17, 1.31315635078607e+17, 1.313156350900132e+17, 1.313156351003258e+17, 1.313156351111071e+17, 1.313156351311071e+17, 1.313156351428257e+17, 1.313156351531383e+17, 1.313156351634508e+17, 1.31315635173607e+17, 1.313156351840758e+17, 1.313156351948571e+17, 1.313156352050132e+17, 1.313156352151695e+17, 1.313156352256383e+17, 1.313156352356383e+17, 1.31315635246107e+17, 1.313156352564195e+17, 1.313156352679821e+17, 1.313156352782945e+17, 1.313156352897007e+17, 1.31315635299857e+17, 1.313156353103258e+17, 1.313156353209508e+17, 1.313156353314194e+17, 1.313156353425133e+17, 1.313156353528257e+17, 1.313156353634508e+17, 1.313156353742321e+17, 1.313156353850132e+17, 1.313156353959508e+17, 1.313156354075133e+17, 1.313156354179821e+17, 1.313156354281382e+17, 1.313156354390757e+17, 1.313156354495446e+17, 1.313156354595444e+17, 1.31315635469857e+17, 1.313156354801695e+17, 1.313156354907945e+17, 1.313156355009508e+17, 1.313156355114195e+17, 1.313156355215757e+17, 1.313156355315757e+17, 1.313156355418883e+17, 1.313156355522008e+17, 1.313156355632945e+17, 1.313156355737632e+17, 1.313156355848571e+17, 1.313156355951695e+17, 1.31315635605482e+17, 1.313156356165757e+17, 1.313156356268883e+17, 1.313156356368882e+17, 1.313156356476695e+17, 1.31315635657982e+17, 1.31315635668607e+17, 1.31315635679232e+17, 1.313156356901695e+17, 1.313156357006382e+17, 1.313156357120444e+17, 1.31315635722357e+17, 1.313156357326696e+17, 1.31315635742982e+17, 1.313156357532945e+17, 1.313156357637633e+17, 1.313156357742319e+17, 1.313156357843882e+17, 1.313156357950132e+17, 1.31315635806107e+17, 1.31315635816107e+17, 1.313156358264195e+17, 1.313156358370445e+17, 1.313156358472008e+17, 1.313156358578258e+17, 1.313156358681382e+17, 1.31315635879232e+17, 1.313156358897007e+17, 1.31315635899857e+17, 1.313156359103258e+17, 1.313156359207945e+17, 1.313156359311069e+17, 1.31315635941732e+17, 1.313156359520445e+17, 1.313156359622008e+17, 1.31315635972357e+17, 1.313156359828257e+17, 1.313156359931383e+17, 1.313156360034508e+17, 1.313156360137633e+17, 1.313156360245444e+17, 1.313156360356383e+17, 1.313156360459507e+17, 1.313156360562633e+17, 1.313156360668882e+17, 1.313156360773571e+17, 1.313156360881382e+17, 1.313156360982945e+17, 1.313156361095444e+17, 1.313156361197007e+17, 1.313156361301695e+17, 1.31315636150482e+17, 1.313156361643882e+17, 1.313156361756383e+17, 1.313156361956383e+17, 1.31315636206107e+17, 1.313156362173571e+17, 1.313156362276695e+17, 1.313156362381382e+17, 1.313156362501695e+17, 1.313156362611071e+17, 1.313156362718883e+17, 1.313156362820444e+17, 1.313156362925132e+17, 1.313156363032945e+17, 1.313156363139195e+17, 1.313156363248571e+17, 1.313156363356383e+17, 1.31315636346107e+17, 1.31315636356732e+17, 1.313156363673571e+17, 1.313156363781382e+17, 1.313156363886071e+17, 1.313156363989196e+17, 1.313156364090757e+17, 1.313156364201695e+17, 1.313156364307945e+17, 1.313156364415758e+17, 1.313156364525133e+17, 1.313156364626694e+17, 1.313156364732945e+17, 1.313156364843882e+17, 1.313156364951695e+17, 1.313156365059508e+17, 1.31315636516107e+17, 1.313156365270445e+17, 1.313156365372008e+17, 1.313156365475132e+17, 1.313156365578258e+17, 1.313156365681382e+17, 1.313156365782945e+17, 1.31315636588607e+17, 1.313156366001696e+17, 1.313156366101695e+17, 1.313156366206382e+17, 1.313156366318883e+17, 1.313156366426696e+17, 1.313156366626696e+17, 1.313156366734508e+17, 1.313156366839195e+17, 1.313156366947007e+17, 1.313156367051695e+17, 1.313156367164195e+17, 1.31315636726732e+17, 1.313156367370445e+17, 1.313156367481382e+17, 1.313156367592321e+17, 1.31315636769857e+17, 1.31315636780482e+17, 1.313156367906382e+17, 1.313156368015757e+17, 1.313156368125132e+17, 1.313156368232945e+17, 1.313156368339195e+17, 1.313156368448571e+17, 1.313156368553257e+17, 1.313156368659507e+17, 1.31315636876107e+17, 1.313156368864195e+17, 1.313156368968882e+17, 1.313156369068883e+17, 1.313156369172008e+17, 1.313156369272008e+17, 1.313156369373571e+17, 1.313156369476695e+17, 1.313156369576695e+17, 1.313156369681382e+17, 1.313156369789194e+17, 1.31315636989857e+17, 1.313156370003258e+17, 1.313156370115757e+17, 1.313156370225133e+17, 1.313156370326696e+17, 1.31315637043607e+17, 1.313156370537632e+17, 1.313156370639195e+17, 1.313156370740758e+17, 1.313156370840756e+17, 1.313156370942321e+17, 1.313156371045445e+17, 1.313156371151695e+17, 1.313156371253257e+17, 1.313156371362632e+17, 1.313156371465757e+17, 1.313156371568882e+17, 1.313156371672008e+17, 1.313156371778258e+17, 1.31315637187982e+17, 1.31315637198607e+17, 1.313156372101695e+17, 1.31315637220482e+17, 1.313156372311069e+17, 1.31315637241732e+17, 1.313156372526696e+17, 1.313156372637632e+17, 1.313156372740758e+17, 1.313156372843882e+17, 1.31315637294857e+17, 1.313156373056383e+17, 1.313156373167319e+17, 1.313156373272008e+17, 1.313156373375132e+17, 1.313156373476695e+17, 1.313156373581382e+17, 1.313156373682945e+17, 1.313156373789196e+17, 1.31315637389857e+17, 1.31315637400482e+17, 1.313156374109508e+17, 1.313156374211069e+17, 1.313156374314195e+17, 1.313156374420445e+17, 1.313156374528257e+17, 1.313156374628257e+17, 1.313156374732945e+17, 1.313156374839195e+17, 1.313156374947007e+17, 1.313156375051695e+17, 1.31315637515482e+17, 1.31315637526107e+17, 1.313156375362633e+17, 1.31315637546732e+17, 1.313156375572008e+17, 1.313156375673571e+17, 1.31315637577982e+17, 1.313156375882944e+17, 1.313156375984508e+17, 1.313156376086071e+17, 1.313156376189196e+17, 1.313156376290757e+17, 1.31315637639232e+17},
			             {1.31315637639232e+17, 1.313156376500132e+17, 1.313156376615758e+17, 1.313156376722007e+17, 1.31315637682357e+17, 1.313156376926694e+17, 1.313156377034508e+17, 1.31315637713607e+17, 1.313156377237632e+17, 1.313156377347007e+17, 1.313156377451695e+17, 1.313156377557944e+17, 1.31315637766107e+17, 1.313156377776695e+17, 1.313156377881382e+17, 1.313156377984507e+17, 1.313156378093883e+17, 1.313156378211071e+17, 1.31315637831732e+17, 1.313156378428257e+17, 1.313156378528257e+17, 1.31315637863607e+17, 1.313156378742321e+17, 1.313156378843884e+17, 1.313156378956383e+17, 1.313156379062633e+17, 1.313156379164195e+17, 1.313156379275132e+17, 1.313156379379821e+17, 1.31315637948607e+17, 1.31315637959232e+17, 1.313156379701695e+17, 1.313156379801695e+17, 1.313156379903258e+17, 1.313156380007945e+17, 1.313156380114195e+17, 1.313156380215758e+17, 1.313156380322007e+17, 1.31315638042357e+17, 1.313156380531383e+17, 1.313156380639195e+17, 1.313156380742319e+17, 1.313156380843882e+17, 1.313156380951695e+17, 1.313156381056383e+17, 1.31315638116107e+17, 1.313156381264195e+17, 1.31315638136732e+17, 1.313156381473571e+17, 1.313156381576695e+17, 1.313156381679821e+17, 1.31315638177982e+17, 1.313156381893883e+17, 1.313156382000132e+17, 1.313156382103258e+17, 1.31315638220482e+17, 1.313156382309507e+17, 1.313156382415758e+17, 1.313156382522007e+17, 1.31315638262982e+17, 1.313156382740758e+17, 1.313156382843882e+17, 1.313156382943884e+17, 1.31315638304857e+17, 1.313156383153257e+17, 1.313156383264195e+17, 1.31315638337982e+17, 1.313156383490758e+17, 1.31315638359232e+17, 1.313156383695444e+17, 1.313156383895444e+17, 1.313156384007945e+17, 1.313156384112632e+17, 1.313156384214195e+17, 1.313156384320444e+17, 1.313156384422008e+17, 1.313156384525133e+17, 1.313156384626696e+17, 1.313156384732945e+17, 1.313156384840758e+17, 1.313156384943882e+17, 1.313156385056381e+17, 1.313156385157944e+17, 1.31315638526107e+17, 1.313156385365756e+17, 1.313156385472008e+17, 1.313156385576695e+17, 1.31315638569232e+17, 1.313156385795444e+17, 1.313156385900132e+17, 1.313156386007945e+17, 1.31315638611732e+17, 1.31315638622982e+17, 1.313156386331382e+17, 1.31315638643607e+17, 1.313156386539195e+17, 1.313156386640756e+17, 1.313156386745445e+17, 1.313156386862633e+17, 1.313156386970445e+17, 1.313156387075133e+17, 1.313156387193882e+17, 1.313156387300133e+17, 1.31315638740482e+17, 1.313156387511069e+17, 1.313156387612632e+17, 1.31315638771732e+17, 1.313156387820444e+17, 1.313156387936069e+17, 1.313156388043882e+17, 1.313156388143884e+17, 1.313156388245445e+17, 1.31315638834857e+17, 1.313156388454821e+17, 1.313156388562633e+17, 1.313156388681382e+17, 1.313156388782945e+17, 1.313156388890757e+17, 1.313156388997007e+17, 1.313156389097007e+17, 1.313156389197007e+17, 1.313156389303258e+17, 1.313156389409508e+17, 1.313156389509508e+17, 1.31315638961732e+17, 1.313156389723571e+17, 1.313156389826696e+17, 1.313156389928257e+17, 1.313156390039195e+17, 1.313156390140756e+17, 1.313156390243882e+17, 1.313156390347007e+17, 1.31315639045482e+17, 1.313156390568883e+17, 1.313156390670445e+17, 1.313156390773569e+17, 1.313156390878258e+17, 1.313156390995444e+17, 1.31315639109857e+17, 1.313156391201695e+17, 1.313156391306382e+17, 1.313156391414195e+17, 1.313156391522008e+17, 1.31315639162982e+17, 1.313156391731383e+17, 1.313156391843884e+17, 1.313156391950132e+17, 1.313156392059507e+17, 1.31315639216732e+17, 1.313156392273569e+17, 1.313156392379821e+17, 1.313156392487633e+17, 1.313156392589194e+17, 1.31315639269232e+17, 1.313156392793883e+17, 1.313156392897007e+17, 1.313156393000133e+17, 1.313156393111069e+17, 1.31315639321732e+17, 1.313156393322008e+17, 1.313156393426694e+17, 1.313156393534508e+17, 1.313156393645444e+17, 1.31315639374857e+17, 1.31315639385482e+17, 1.31315639396107e+17, 1.313156394064195e+17, 1.313156394172008e+17, 1.313156394275133e+17, 1.313156394387633e+17, 1.313156394489196e+17, 1.313156394597007e+17, 1.313156394703258e+17, 1.313156394812632e+17, 1.31315639491732e+17, 1.313156395022008e+17, 1.313156395126696e+17, 1.313156395228257e+17, 1.313156395328257e+17, 1.313156395428257e+17, 1.313156395628257e+17, 1.313156395747008e+17, 1.313156395856383e+17, 1.313156395962633e+17, 1.313156396065757e+17, 1.313156396165757e+17, 1.31315639626732e+17, 1.313156396368882e+17, 1.313156396473571e+17, 1.313156396576695e+17, 1.313156396681382e+17, 1.313156396790757e+17, 1.313156396897007e+17, 1.313156397006382e+17, 1.313156397107945e+17, 1.313156397209508e+17, 1.313156397317321e+17, 1.313156397428257e+17, 1.313156397531383e+17, 1.313156397634508e+17, 1.313156397739195e+17, 1.31315639784857e+17, 1.31315639795482e+17, 1.313156398065757e+17, 1.313156398172008e+17, 1.313156398273571e+17, 1.313156398375133e+17, 1.313156398476695e+17, 1.313156398589196e+17, 1.31315639869232e+17, 1.313156398793883e+17, 1.313156398903258e+17, 1.313156399014195e+17, 1.313156399115758e+17, 1.313156399225133e+17, 1.313156399328259e+17, 1.313156399431383e+17, 1.313156399534508e+17, 1.313156399642319e+17, 1.313156399745445e+17, 1.313156399850132e+17, 1.313156399959507e+17, 1.31315640006107e+17, 1.313156400162633e+17, 1.313156400262632e+17, 1.313156400368882e+17, 1.313156400472008e+17, 1.313156400578257e+17, 1.313156400682945e+17, 1.313156400795444e+17, 1.31315640089857e+17, 1.313156401003258e+17, 1.313156401112632e+17, 1.313156401222007e+17, 1.313156401325133e+17, 1.31315640142982e+17, 1.313156401531382e+17, 1.313156401637633e+17, 1.313156401740758e+17, 1.313156401842319e+17, 1.313156401943882e+17, 1.313156402057946e+17, 1.31315640216107e+17, 1.313156402265757e+17, 1.313156402382945e+17, 1.313156402484507e+17, 1.313156402589194e+17, 1.313156402690757e+17, 1.31315640279232e+17, 1.313156402895444e+17, 1.313156403007944e+17, 1.313156403115757e+17, 1.313156403218883e+17, 1.31315640332357e+17, 1.313156403437632e+17, 1.313156403539195e+17, 1.313156403640758e+17, 1.313156403742319e+17, 1.313156403843882e+17, 1.313156403947008e+17, 1.313156404050132e+17, 1.313156404153257e+17, 1.31315640426107e+17, 1.313156404368882e+17, 1.313156404478257e+17, 1.31315640457982e+17, 1.313156404682944e+17, 1.313156404789196e+17, 1.313156404895444e+17, 1.313156405001695e+17, 1.313156405103258e+17, 1.313156405206382e+17, 1.313156405309507e+17, 1.313156405409508e+17, 1.313156405515757e+17, 1.313156405620444e+17, 1.31315640572357e+17, 1.313156405828257e+17, 1.313156405939195e+17, 1.313156406042321e+17, 1.313156406143882e+17, 1.313156406245444e+17, 1.31315640634857e+17, 1.313156406451695e+17, 1.313156406556383e+17, 1.313156406659507e+17, 1.313156406764196e+17, 1.31315640686732e+17, 1.313156406968882e+17, 1.313156407078257e+17, 1.31315640719232e+17, 1.313156407297007e+17, 1.31315640739857e+17, 1.313156407503256e+17, 1.313156407614195e+17, 1.31315640772357e+17, 1.31315640782982e+17, 1.313156407934508e+17, 1.313156408037632e+17, 1.313156408140756e+17, 1.313156408245445e+17, 1.31315640834857e+17, 1.31315640845482e+17, 1.313156408564195e+17, 1.313156408672008e+17, 1.313156408773569e+17, 1.313156408889194e+17, 1.31315640899232e+17, 1.313156409095444e+17, 1.313156409200133e+17, 1.313156409317321e+17, 1.31315640942982e+17, 1.313156409531383e+17, 1.313156409647007e+17, 1.313156409753258e+17, 1.313156409859507e+17, 1.313156409964195e+17, 1.313156410065757e+17, 1.313156410168883e+17, 1.313156410275133e+17, 1.313156410381382e+17, 1.313156410489196e+17, 1.313156410620444e+17, 1.313156410726696e+17, 1.31315641083607e+17, 1.313156410937633e+17, 1.313156411040758e+17, 1.313156411147007e+17, 1.31315641124857e+17, 1.313156411351695e+17, 1.313156411457944e+17, 1.313156411570445e+17, 1.313156411679821e+17, 1.313156411782945e+17, 1.313156411884507e+17, 1.31315641198607e+17, 1.313156412097007e+17, 1.313156412201695e+17, 1.313156412306383e+17, 1.31315641241732e+17, 1.313156412518883e+17, 1.31315641262357e+17, 1.313156412725133e+17, 1.313156412826696e+17, 1.313156412928257e+17, 1.313156413028257e+17, 1.31315641312982e+17, 1.313156413231383e+17, 1.313156413336069e+17, 1.313156413439195e+17, 1.313156413543884e+17, 1.313156413650132e+17, 1.313156413764195e+17, 1.313156413868883e+17, 1.313156413970445e+17, 1.313156414075132e+17, 1.313156414178258e+17, 1.313156414287633e+17, 1.313156414395444e+17, 1.313156414497007e+17, 1.313156414600133e+17, 1.313156414701695e+17, 1.313156414806382e+17, 1.313156414909507e+17, 1.313156415022007e+17, 1.31315641512357e+17, 1.313156415226696e+17, 1.313156415334508e+17, 1.313156415445445e+17, 1.313156415553257e+17, 1.313156415665757e+17, 1.31315641576732e+17, 1.313156415870446e+17, 1.313156415976695e+17, 1.313156416078258e+17, 1.313156416182944e+17, 1.31315641628607e+17, 1.313156416387633e+17, 1.313156416495444e+17, 1.31315641659857e+17, 1.313156416700133e+17, 1.313156416806383e+17, 1.313156416918883e+17, 1.313156417026696e+17, 1.313156417132945e+17, 1.313156417236069e+17, 1.313156417340758e+17, 1.313156417442319e+17, 1.313156417547008e+17, 1.313156417653257e+17, 1.313156417765757e+17, 1.313156417870445e+17, 1.313156417976695e+17, 1.313156418084507e+17, 1.31315641818607e+17, 1.313156418293883e+17, 1.313156418400132e+17, 1.313156418509508e+17, 1.313156418620444e+17, 1.313156418720445e+17, 1.31315641882357e+17, 1.313156418925132e+17, 1.313156419028257e+17, 1.313156419137632e+17, 1.313156419248571e+17, 1.313156419350132e+17, 1.313156419459507e+17, 1.313156419570446e+17, 1.313156419672008e+17, 1.31315641977982e+17, 1.31315641989232e+17, 1.313156419995446e+17, 1.31315642009857e+17, 1.313156420204819e+17, 1.313156420311071e+17, 1.313156420425132e+17, 1.313156420528257e+17, 1.313156420631382e+17, 1.313156420734508e+17, 1.31315642083607e+17, 1.313156420947008e+17, 1.31315642106107e+17, 1.313156421164195e+17, 1.313156421273571e+17, 1.313156421375133e+17, 1.313156421476695e+17, 1.313156421584507e+17, 1.31315642169232e+17, 1.313156421804819e+17, 1.313156421911071e+17, 1.313156422014195e+17, 1.313156422126694e+17, 1.31315642222982e+17, 1.313156422334508e+17, 1.31315642243607e+17, 1.313156422539195e+17, 1.313156422642319e+17, 1.313156422742321e+17, 1.313156422847008e+17, 1.313156422951694e+17, 1.31315642305482e+17, 1.313156423157944e+17, 1.313156423264196e+17, 1.313156423373571e+17, 1.313156423478258e+17, 1.313156423584507e+17, 1.313156423690757e+17, 1.31315642379857e+17, 1.313156423901696e+17, 1.31315642400482e+17, 1.313156424107945e+17, 1.313156424209507e+17, 1.313156424314195e+17, 1.313156424425133e+17, 1.313156424528257e+17, 1.313156424631383e+17, 1.313156424734508e+17, 1.313156424934508e+17, 1.313156425037633e+17, 1.313156425142321e+17, 1.313156425342321e+17, 1.313156425445445e+17, 1.313156425547007e+17, 1.313156425650132e+17, 1.313156425764195e+17, 1.313156425872008e+17, 1.313156425984507e+17, 1.313156426090757e+17, 1.313156426193883e+17, 1.313156426293883e+17, 1.313156426406383e+17, 1.313156426514195e+17, 1.313156426628257e+17, 1.31315642672982e+17, 1.313156426847007e+17, 1.31315642694857e+17, 1.313156427050132e+17, 1.313156427151695e+17, 1.313156427257944e+17, 1.31315642736107e+17, 1.313156427462633e+17, 1.313156427565757e+17, 1.313156427670445e+17, 1.313156427775132e+17, 1.31315642787982e+17, 1.313156427981382e+17, 1.31315642808607e+17, 1.313156428193883e+17, 1.313156428301696e+17, 1.313156428406382e+17, 1.313156428514195e+17, 1.313156428618883e+17, 1.31315642872357e+17, 1.313156428828257e+17, 1.313156428936069e+17, 1.313156429037632e+17, 1.313156429139195e+17, 1.313156429251694e+17, 1.313156429353257e+17, 1.313156429457944e+17, 1.313156429564196e+17, 1.313156429673571e+17, 1.313156429778258e+17, 1.313156429881382e+17, 1.31315642999232e+17, 1.313156430106383e+17, 1.31315643021732e+17, 1.31315643032357e+17, 1.313156430426696e+17, 1.313156430531383e+17, 1.313156430634508e+17, 1.313156430737633e+17, 1.313156430842319e+17, 1.313156430943882e+17, 1.313156431047008e+17, 1.313156431150132e+17, 1.313156431257946e+17, 1.313156431370445e+17, 1.313156431473571e+17, 1.313156431576695e+17, 1.313156431684508e+17, 1.31315643178607e+17, 1.313156431889194e+17, 1.313156431995446e+17, 1.313156432103258e+17, 1.313156432204819e+17, 1.313156432311071e+17, 1.313156432414195e+17, 1.313156432515758e+17, 1.313156432618883e+17, 1.313156432731382e+17, 1.313156432839195e+17, 1.313156432940758e+17, 1.313156433050132e+17, 1.313156433150132e+17, 1.313156433256383e+17, 1.313156433370445e+17, 1.313156433475132e+17, 1.313156433576695e+17, 1.313156433678258e+17, 1.313156433779821e+17, 1.313156433884508e+17, 1.313156433987633e+17, 1.313156434097007e+17, 1.313156434203256e+17, 1.313156434307945e+17, 1.31315643441732e+17, 1.313156434518883e+17, 1.31315643462357e+17, 1.313156434726694e+17, 1.31315643482982e+17, 1.313156434937632e+17, 1.313156435042319e+17, 1.313156435147008e+17, 1.313156435265757e+17, 1.313156435372008e+17, 1.313156435481384e+17, 1.313156435582944e+17, 1.313156435684508e+17, 1.313156435790758e+17, 1.313156435893883e+17, 1.313156435997007e+17, 1.313156436100133e+17, 1.313156436203258e+17, 1.313156436306382e+17, 1.313156436418883e+17, 1.313156436522007e+17, 1.313156436626694e+17, 1.313156436731382e+17, 1.313156436832945e+17, 1.313156436934508e+17, 1.31315643703607e+17, 1.313156437137632e+17, 1.313156437240756e+17, 1.313156437351695e+17, 1.31315643745482e+17, 1.31315643756107e+17, 1.313156437675133e+17, 1.313156437781382e+17, 1.313156437893883e+17, 1.313156437997007e+17, 1.313156438101695e+17, 1.31315643820482e+17, 1.313156438312634e+17, 1.313156438415758e+17, 1.31315643851732e+17, 1.31315643862982e+17, 1.31315643873607e+17, 1.313156438837632e+17, 1.313156438940756e+17, 1.313156439051694e+17, 1.313156439157946e+17, 1.313156439264195e+17, 1.31315643936732e+17, 1.313156439468883e+17, 1.313156439573569e+17, 1.313156439679821e+17, 1.313156439784508e+17, 1.313156439890757e+17, 1.31315643999857e+17, 1.31315644010482e+17, 1.313156440212632e+17, 1.313156440315757e+17, 1.313156440425133e+17, 1.313156440526694e+17, 1.313156440632945e+17, 1.313156440734508e+17, 1.313156440836069e+17, 1.313156440942321e+17, 1.31315644104857e+17, 1.31315644115482e+17, 1.31315644126107e+17, 1.313156441370445e+17, 1.313156441475132e+17, 1.313156441576695e+17, 1.313156441687633e+17, 1.313156441790757e+17, 1.31315644189857e+17, 1.313156442000133e+17, 1.313156442114195e+17, 1.313156442228257e+17, 1.313156442340758e+17, 1.313156442442321e+17, 1.313156442545445e+17, 1.31315644264857e+17, 1.313156442750132e+17, 1.31315644285482e+17, 1.313156442956383e+17, 1.31315644306107e+17, 1.313156443165757e+17, 1.313156443268883e+17, 1.313156443376695e+17, 1.313156443481382e+17, 1.313156443582944e+17, 1.313156443684507e+17, 1.313156443793883e+17, 1.313156443903258e+17, 1.313156444007945e+17, 1.313156444111069e+17, 1.313156444212632e+17, 1.313156444318883e+17, 1.313156444422007e+17, 1.31315644452357e+17, 1.313156444625133e+17, 1.31315644472982e+17, 1.313156444832945e+17, 1.31315644493607e+17, 1.313156445042321e+17, 1.313156445147008e+17, 1.313156445264195e+17, 1.313156445372008e+17, 1.313156445478257e+17, 1.313156445589196e+17, 1.31315644569232e+17, 1.313156445795444e+17, 1.313156445897007e+17, 1.313156446000133e+17, 1.313156446101696e+17, 1.31315644620482e+17, 1.313156446309508e+17, 1.313156446415758e+17, 1.313156446522007e+17, 1.31315644662982e+17, 1.313156446736069e+17, 1.313156446942319e+17, 1.313156447043882e+17, 1.313156447145445e+17, 1.313156447247007e+17, 1.313156447351695e+17, 1.313156447457944e+17, 1.313156447564196e+17, 1.313156447665756e+17, 1.313156447778258e+17, 1.313156447879821e+17, 1.313156447990757e+17, 1.31315644809232e+17, 1.31315644819857e+17, 1.313156448312634e+17, 1.31315644841732e+17, 1.31315644852357e+17, 1.313156448625132e+17, 1.31315644873607e+17, 1.313156448840758e+17, 1.313156448943884e+17, 1.313156449047008e+17, 1.313156449151695e+17, 1.313156449257944e+17, 1.313156449364195e+17, 1.31315644946732e+17, 1.313156449570445e+17, 1.313156449673571e+17, 1.31315644977982e+17, 1.313156449881382e+17, 1.313156449984507e+17, 1.313156450087633e+17, 1.313156450189196e+17, 1.313156450293883e+17, 1.313156450397007e+17, 1.313156450500133e+17, 1.313156450601696e+17, 1.313156450706382e+17, 1.313156450807945e+17, 1.313156450915757e+17, 1.313156451026696e+17, 1.313156451134508e+17, 1.313156451237632e+17, 1.313156451340758e+17, 1.313156451443882e+17, 1.313156451550132e+17, 1.313156451656383e+17, 1.313156451759507e+17, 1.313156451872008e+17, 1.313156451984507e+17, 1.31315645208607e+17, 1.313156452189196e+17, 1.313156452290757e+17, 1.313156452393883e+17, 1.313156452497007e+17, 1.31315645259857e+17, 1.313156452703258e+17, 1.313156452806382e+17, 1.313156452907945e+17, 1.313156453015758e+17, 1.313156453118883e+17, 1.313156453225133e+17, 1.313156453337633e+17, 1.313156453440758e+17, 1.313156453547007e+17, 1.313156453650132e+17, 1.313156453756383e+17, 1.313156453856383e+17, 1.313156453962633e+17, 1.313156454068882e+17, 1.313156454176695e+17, 1.31315645427982e+17, 1.313156454381382e+17, 1.313156454481382e+17, 1.313156454587633e+17, 1.313156454690758e+17, 1.313156454797007e+17, 1.313156454909508e+17, 1.313156455012634e+17, 1.313156455114195e+17, 1.313156455215757e+17, 1.313156455325133e+17, 1.313156455426696e+17, 1.313156455532945e+17, 1.313156455637633e+17, 1.313156455745445e+17, 1.313156455847008e+17, 1.313156455950132e+17, 1.313156456050132e+17, 1.31315645615482e+17, 1.313156456267319e+17, 1.313156456373571e+17, 1.313156456489196e+17, 1.313156456601695e+17, 1.313156456703258e+17, 1.31315645680482e+17, 1.313156456911069e+17, 1.313156457015757e+17, 1.31315645711732e+17, 1.313156457226694e+17, 1.313156457331382e+17, 1.313156457432945e+17, 1.313156457540758e+17, 1.313156457642321e+17, 1.313156457750132e+17, 1.313156457859507e+17, 1.313156457962633e+17, 1.313156458065757e+17, 1.313156458176695e+17, 1.31315645827982e+17, 1.313156458381382e+17, 1.313156458482945e+17, 1.313156458584508e+17, 1.31315645869232e+17, 1.313156458795444e+17, 1.313156458897007e+17, 1.313156459000133e+17, 1.313156459109508e+17, 1.313156459212632e+17, 1.313156459312632e+17, 1.313156459418883e+17, 1.313156459522007e+17, 1.313156459626694e+17, 1.313156459731382e+17, 1.313156459832945e+17, 1.313156459934508e+17, 1.313156460037633e+17, 1.313156460142319e+17, 1.313156460245445e+17, 1.313156460350132e+17, 1.313156460450132e+17, 1.313156460564195e+17, 1.313156460672008e+17, 1.313156460776695e+17, 1.313156460884507e+17, 1.31315646099232e+17, 1.313156461093883e+17, 1.313156461197007e+17, 1.313156461300133e+17, 1.313156461401695e+17, 1.313156461504819e+17, 1.313156461606382e+17, 1.313156461714195e+17, 1.313156461815758e+17, 1.31315646192357e+17, 1.31315646202982e+17, 1.313156462140758e+17, 1.313156462242321e+17, 1.313156462345445e+17, 1.313156462445445e+17, 1.313156462545445e+17, 1.313156462647007e+17, 1.313156462750132e+17, 1.313156462851695e+17, 1.313156462956381e+17, 1.313156463057944e+17, 1.313156463164195e+17, 1.313156463265757e+17, 1.313156463365757e+17, 1.313156463470445e+17, 1.313156463572008e+17, 1.313156463681384e+17, 1.31315646378607e+17, 1.313156463887633e+17, 1.31315646399232e+17, 1.31315646409857e+17, 1.313156464203258e+17, 1.313156464304819e+17, 1.313156464411071e+17, 1.313156464512632e+17, 1.313156464614195e+17, 1.31315646471732e+17, 1.313156464822007e+17, 1.313156464926696e+17, 1.313156465039195e+17, 1.313156465140758e+17, 1.313156465243884e+17, 1.313156465347008e+17, 1.31315646544857e+17, 1.31315646555482e+17, 1.313156465668883e+17, 1.313156465775132e+17, 1.313156465878257e+17, 1.31315646597982e+17, 1.313156466084507e+17, 1.313156466187633e+17, 1.313156466293883e+17, 1.313156466400133e+17, 1.313156466503258e+17, 1.31315646660482e+17, 1.313156466707945e+17, 1.313156466814194e+17, 1.313156466914195e+17, 1.313156467020444e+17, 1.313156467131383e+17, 1.313156467237632e+17, 1.313156467340758e+17, 1.313156467442321e+17, 1.313156467545445e+17, 1.313156467647007e+17, 1.313156467751695e+17, 1.313156467853257e+17, 1.313156467957946e+17, 1.313156468078257e+17, 1.313156468178258e+17, 1.313156468279821e+17, 1.313156468389196e+17, 1.313156468490757e+17, 1.31315646859232e+17, 1.313156468700133e+17, 1.313156468801695e+17, 1.313156468903258e+17, 1.313156469015758e+17, 1.313156469122007e+17, 1.313156469228257e+17, 1.31315646932982e+17, 1.31315646943607e+17, 1.313156469540758e+17, 1.313156469642321e+17, 1.313156469747007e+17, 1.313156469857944e+17, 1.313156469959507e+17, 1.313156470065757e+17, 1.31315647016732e+17, 1.31315647026732e+17, 1.313156470370445e+17, 1.313156470482945e+17, 1.31315647058607e+17, 1.313156470689194e+17, 1.313156470793882e+17, 1.313156470900133e+17, 1.313156471001696e+17, 1.313156471103258e+17, 1.31315647120482e+17, 1.313156471307945e+17, 1.313156471412632e+17, 1.313156471515757e+17, 1.313156471625132e+17, 1.313156471732945e+17, 1.31315647183607e+17, 1.313156471940756e+17, 1.313156472042321e+17, 1.313156472147008e+17, 1.313156472251694e+17, 1.313156472357944e+17, 1.313156472465757e+17, 1.313156472567319e+17, 1.313156472670445e+17, 1.313156472773569e+17, 1.313156472879821e+17, 1.313156472987633e+17, 1.313156473095444e+17, 1.313156473203258e+17, 1.313156473311071e+17, 1.31315647341732e+17, 1.313156473523571e+17, 1.313156473626696e+17, 1.313156473726694e+17, 1.313156473832946e+17, 1.313156473937632e+17, 1.313156474042321e+17, 1.313156474143884e+17, 1.31315647424857e+17, 1.31315647436107e+17, 1.313156474464196e+17, 1.31315647456732e+17, 1.313156474672008e+17, 1.31315647477982e+17, 1.313156474882945e+17, 1.313156474984507e+17, 1.31315647508607e+17, 1.313156475187633e+17, 1.313156475290757e+17, 1.313156475398569e+17, 1.313156475503258e+17, 1.313156475609508e+17, 1.313156475717321e+17, 1.313156475820445e+17, 1.313156475926694e+17, 1.313156476028257e+17, 1.313156476132945e+17, 1.313156476237632e+17, 1.313156476340758e+17, 1.313156476447008e+17, 1.313156476550132e+17, 1.313156476653258e+17, 1.313156476756383e+17, 1.31315647686107e+17, 1.313156476972006e+17, 1.313156477078258e+17, 1.313156477178257e+17, 1.313156477284508e+17, 1.313156477389194e+17, 1.313156477495446e+17, 1.313156477597007e+17, 1.313156477701695e+17, 1.313156477812632e+17, 1.313156477915758e+17, 1.31315647802357e+17, 1.313156478128257e+17, 1.313156478234508e+17, 1.313156478337632e+17, 1.313156478450132e+17, 1.313156478553258e+17, 1.31315647865482e+17, 1.313156478756383e+17, 1.313156478859507e+17, 1.313156478968882e+17, 1.313156479078258e+17, 1.313156479182944e+17, 1.313156479284507e+17, 1.313156479387633e+17, 1.313156479489196e+17, 1.313156479590757e+17, 1.313156479695444e+17, 1.313156479797007e+17, 1.313156479900132e+17, 1.313156480007945e+17, 1.313156480111071e+17, 1.313156480217321e+17, 1.31315648031732e+17, 1.313156480425133e+17, 1.31315648052982e+17, 1.313156480634508e+17, 1.31315648073607e+17, 1.313156480842319e+17, 1.313156480943882e+17, 1.313156481047008e+17, 1.313156481151694e+17, 1.313156481259507e+17, 1.31315648136107e+17, 1.313156481464196e+17, 1.313156481568882e+17, 1.313156481681382e+17, 1.313156481781382e+17, 1.313156481890757e+17, 1.313156481997007e+17, 1.313156482104819e+17, 1.313156482214195e+17, 1.313156482322008e+17, 1.313156482423571e+17, 1.313156482526696e+17, 1.313156482631383e+17, 1.313156482740758e+17, 1.313156482842321e+17, 1.313156482947008e+17, 1.313156483051695e+17, 1.313156483151695e+17, 1.31315648326107e+17, 1.313156483375132e+17, 1.313156483475132e+17, 1.313156483578258e+17, 1.313156483687633e+17, 1.31315648379857e+17, 1.313156483901695e+17, 1.313156484009508e+17, 1.313156484112632e+17, 1.313156484214195e+17, 1.313156484318883e+17, 1.313156484422008e+17, 1.313156484525133e+17, 1.313156484628259e+17, 1.313156484732945e+17, 1.313156484843882e+17, 1.313156484947007e+17, 1.313156485050132e+17, 1.313156485162633e+17, 1.313156485264195e+17, 1.31315648536732e+17, 1.313156485470445e+17, 1.313156485573569e+17, 1.313156485676695e+17, 1.31315648578607e+17, 1.313156485887633e+17, 1.313156485995444e+17, 1.313156486100133e+17, 1.313156486203258e+17, 1.313156486312632e+17, 1.313156486414195e+17, 1.313156486515757e+17, 1.313156486625133e+17, 1.313156486728257e+17, 1.313156486828257e+17, 1.313156486931383e+17, 1.31315648703607e+17, 1.313156487142319e+17, 1.313156487243882e+17, 1.313156487347008e+17, 1.313156487450132e+17, 1.31315648756732e+17, 1.313156487673571e+17, 1.313156487776695e+17, 1.313156487881382e+17, 1.313156487987633e+17, 1.313156488090758e+17, 1.313156488197007e+17, 1.31315648830482e+17, 1.313156488412632e+17, 1.31315648851732e+17, 1.31315648861732e+17, 1.313156488720444e+17, 1.313156488828257e+17, 1.31315648892982e+17, 1.313156489031382e+17, 1.313156489134508e+17, 1.31315648923607e+17, 1.313156489340756e+17, 1.313156489450132e+17, 1.31315648955482e+17, 1.313156489659508e+17, 1.313156489765757e+17, 1.313156489868882e+17, 1.313156489972008e+17, 1.31315649007982e+17, 1.313156490182945e+17, 1.313156490284508e+17, 1.313156490390757e+17, 1.313156490501695e+17, 1.313156490604819e+17, 1.313156490711069e+17, 1.313156490812632e+17, 1.313156490922008e+17, 1.31315649102982e+17, 1.313156491132945e+17, 1.313156491236069e+17, 1.313156491337632e+17, 1.313156491442319e+17, 1.313156491547008e+17, 1.313156491650132e+17, 1.31315649175482e+17, 1.313156491864196e+17, 1.313156491975132e+17, 1.313156492076695e+17, 1.313156492182944e+17, 1.31315649229232e+17, 1.313156492395444e+17, 1.313156492493882e+17, 1.313156492603258e+17, 1.31315649270482e+17, 1.31315649280482e+17, 1.313156492903258e+17, 1.313156493003258e+17, 1.313156493103258e+17, 1.31315649321732e+17, 1.31315649332357e+17, 1.313156493432945e+17, 1.31315649353607e+17, 1.313156493639195e+17, 1.313156493739195e+17, 1.313156493836069e+17, 1.313156493931383e+17, 1.31315649402357e+17, 1.313156494120445e+17, 1.313156494218883e+17, 1.313156494307945e+17, 1.313156494409508e+17, 1.313156494500133e+17, 1.313156494595444e+17, 1.313156494687633e+17, 1.313156494779821e+17, 1.31315649487982e+17, 1.313156494981382e+17, 1.31315649509232e+17, 1.313156495181382e+17, 1.313156495275132e+17, 1.313156495368883e+17, 1.313156495468883e+17, 1.313156495562633e+17, 1.313156495657944e+17, 1.313156495751695e+17, 1.313156495847007e+17, 1.31315649593607e+17, 1.313156496039195e+17, 1.313156496132945e+17, 1.31315649622357e+17, 1.313156496318883e+17, 1.313156496409508e+17, 1.313156496501695e+17, 1.313156496593882e+17, 1.313156496695444e+17, 1.313156496789194e+17, 1.313156496882945e+17, 1.313156496978258e+17, 1.31315649707982e+17, 1.313156497195444e+17, 1.313156497300133e+17, 1.313156497412632e+17, 1.31315649751732e+17, 1.313156497620444e+17, 1.313156497726696e+17, 1.313156497839195e+17, 1.313156497942319e+17, 1.313156498051695e+17, 1.313156498157946e+17, 1.313156498265757e+17, 1.313156498372008e+17, 1.313156498484507e+17, 1.313156498590757e+17, 1.31315649870482e+17, 1.313156498815757e+17, 1.313156498922007e+17, 1.313156499036069e+17, 1.313156499153258e+17, 1.313156499262633e+17, 1.313156499370445e+17, 1.313156499476695e+17, 1.313156499582944e+17, 1.313156499690757e+17, 1.31315649980482e+17, 1.313156499911069e+17, 1.313156500022008e+17, 1.313156500134508e+17, 1.31315650024857e+17, 1.313156500356383e+17, 1.313156500464195e+17, 1.313156500570445e+17, 1.313156500676695e+17, 1.313156500778257e+17, 1.313156500881382e+17, 1.313156500982945e+17, 1.313156501086071e+17, 1.313156501190757e+17, 1.313156501306383e+17, 1.313156501414195e+17, 1.313156501515757e+17, 1.31315650161732e+17, 1.313156501718883e+17, 1.31315650182357e+17, 1.313156501926696e+17, 1.31315650203607e+17, 1.313156502139195e+17, 1.313156502245445e+17, 1.313156502347007e+17, 1.313156502456383e+17, 1.313156502564195e+17, 1.313156502668882e+17, 1.31315650277982e+17, 1.313156502893882e+17, 1.313156503012632e+17, 1.313156503132946e+17, 1.313156503256383e+17, 1.313156503384507e+17, 1.313156503512632e+17, 1.313156503639195e+17, 1.313156503762632e+17, 1.313156503882945e+17, 1.313156504004819e+17, 1.313156504125133e+17, 1.313156504245445e+17, 1.313156504368883e+17, 1.31315650449232e+17, 1.313156504618883e+17, 1.313156504739195e+17, 1.31315650486107e+17, 1.313156504982945e+17, 1.313156505106382e+17, 1.313156505228257e+17, 1.31315650534857e+17, 1.313156505473571e+17, 1.313156505593883e+17, 1.313156505715758e+17, 1.31315650583607e+17, 1.313156505962632e+17, 1.313156506089196e+17, 1.313156506211069e+17, 1.313156506332945e+17, 1.313156506453257e+17, 1.313156506573571e+17, 1.313156506693883e+17, 1.313156506814195e+17, 1.313156506934508e+17, 1.31315650705482e+17, 1.313156507184508e+17, 1.313156507312634e+17, 1.31315650743607e+17, 1.313156507559507e+17, 1.31315650767982e+17, 1.313156507801695e+17, 1.31315650792357e+17, 1.313156508045445e+17, 1.313156508168883e+17, 1.313156508290757e+17, 1.313156508412634e+17, 1.313156508532945e+17, 1.31315650865482e+17, 1.313156508778258e+17, 1.313156508903258e+17, 1.313156509025133e+17, 1.313156509145445e+17, 1.313156509268883e+17, 1.313156509389196e+17, 1.313156509514195e+17, 1.313156509639195e+17, 1.31315650976107e+17, 1.313156509881382e+17, 1.313156510007945e+17, 1.313156510129819e+17, 1.313156510251695e+17, 1.313156510375133e+17, 1.313156510495446e+17, 1.313156510620444e+17, 1.313156510742319e+17, 1.31315651086732e+17, 1.313156510990757e+17, 1.313156511114195e+17, 1.31315651123607e+17, 1.313156511356383e+17, 1.313156511481382e+17, 1.31315651160482e+17, 1.313156511726694e+17, 1.31315651184857e+17, 1.313156511972008e+17, 1.313156512093883e+17, 1.31315651221732e+17, 1.313156512343884e+17, 1.313156512465757e+17, 1.313156512587633e+17, 1.313156512711069e+17, 1.313156512834508e+17, 1.31315651295482e+17, 1.313156513078258e+17, 1.31315651320482e+17, 1.31315651332982e+17, 1.313156513451694e+17, 1.313156513575132e+17, 1.31315651369857e+17, 1.313156513820445e+17, 1.313156513940758e+17, 1.313156514064196e+17, 1.313156514189196e+17, 1.313156514309507e+17, 1.313156514432945e+17, 1.313156514559507e+17, 1.31315651467982e+17, 1.313156514803258e+17, 1.31315651492357e+17, 1.313156515043882e+17, 1.31315651516732e+17, 1.313156515287633e+17, 1.313156515409508e+17, 1.31315651552982e+17, 1.313156515650132e+17, 1.313156515772008e+17, 1.313156515900132e+17, 1.313156516020445e+17, 1.313156516147008e+17, 1.31315651626732e+17, 1.313156516387633e+17, 1.313156516507945e+17, 1.313156516628257e+17, 1.313156516748571e+17, 1.313156516872008e+17, 1.313156516995444e+17, 1.313156517117321e+17, 1.313156517242319e+17, 1.313156517362633e+17, 1.313156517487633e+17, 1.313156517607944e+17, 1.313156517732945e+17, 1.313156517853258e+17, 1.313156517973571e+17, 1.313156518095446e+17, 1.313156518218883e+17, 1.313156518340758e+17, 1.31315651846107e+17, 1.313156518582945e+17, 1.313156518703258e+17, 1.313156518826694e+17, 1.31315651894857e+17, 1.313156519068883e+17, 1.313156519193882e+17, 1.313156519320444e+17, 1.31315651944857e+17, 1.313156519568883e+17, 1.313156519693883e+17, 1.313156519815758e+17, 1.31315651993607e+17, 1.313156520059508e+17, 1.313156520179821e+17, 1.313156520301696e+17, 1.31315652042357e+17, 1.313156520543884e+17, 1.313156520665757e+17, 1.313156520790757e+17, 1.313156520912632e+17, 1.313156521034508e+17, 1.31315652115482e+17, 1.313156521275132e+17, 1.313156521397007e+17, 1.313156521518883e+17, 1.313156521639195e+17, 1.31315652176107e+17, 1.313156521884507e+17, 1.31315652200482e+17, 1.313156522125133e+17, 1.31315652224857e+17, 1.313156522368882e+17, 1.31315652249232e+17, 1.313156522615758e+17, 1.313156522739195e+17, 1.313156522859507e+17, 1.313156522979821e+17, 1.313156523103258e+17, 1.313156523223571e+17, 1.313156523347008e+17, 1.31315652346732e+17, 1.313156523590757e+17, 1.313156523714195e+17, 1.313156523837633e+17, 1.313156523957946e+17, 1.313156524079821e+17, 1.313156524201695e+17, 1.31315652432357e+17, 1.313156524445445e+17, 1.313156524565757e+17, 1.31315652468607e+17, 1.313156524807945e+17, 1.313156524931383e+17, 1.313156525057946e+17, 1.313156525179821e+17, 1.31315652530482e+17, 1.313156525425133e+17, 1.313156525545445e+17, 1.31315652566732e+17, 1.313156525789196e+17, 1.313156525914195e+17, 1.31315652603607e+17, 1.313156526157946e+17, 1.313156526281382e+17, 1.313156526403258e+17, 1.31315652652357e+17, 1.313156526647008e+17, 1.31315652676732e+17, 1.313156526887633e+17, 1.313156527009508e+17, 1.313156527134508e+17, 1.313156527256383e+17, 1.313156527378258e+17, 1.313156527503258e+17, 1.31315652762357e+17, 1.313156527743882e+17, 1.313156527865757e+17, 1.313156527987633e+17, 1.313156528109508e+17, 1.31315652822982e+17, 1.313156528353257e+17, 1.313156528475132e+17, 1.313156528597007e+17, 1.31315652871732e+17, 1.313156528837632e+17, 1.313156528962632e+17, 1.31315652908607e+17, 1.313156529207945e+17, 1.313156529328257e+17, 1.31315652945482e+17, 1.313156529575132e+17, 1.313156529697007e+17, 1.31315652981732e+17, 1.313156529937632e+17, 1.31315653006107e+17, 1.313156530187633e+17, 1.313156530307945e+17, 1.313156530426694e+17, 1.313156530547007e+17, 1.31315653066732e+17, 1.313156530787633e+17, 1.313156530907945e+17, 1.313156531028257e+17},
			             {1.31315637639232e+17, 1.313156376500132e+17, 1.313156376615758e+17, 1.313156376722007e+17, 1.31315637682357e+17, 1.313156376926694e+17, 1.313156377034508e+17, 1.31315637713607e+17, 1.313156377237632e+17, 1.313156377347007e+17, 1.313156377451695e+17, 1.313156377557944e+17, 1.31315637766107e+17, 1.313156377776695e+17, 1.313156377881382e+17, 1.313156377984507e+17, 1.313156378093883e+17, 1.313156378211071e+17, 1.31315637831732e+17, 1.313156378428257e+17, 1.313156378528257e+17, 1.31315637863607e+17, 1.313156378742321e+17, 1.313156378843884e+17, 1.313156378956383e+17, 1.313156379062633e+17, 1.313156379164195e+17, 1.313156379275132e+17, 1.313156379379821e+17, 1.31315637948607e+17, 1.31315637959232e+17, 1.313156379701695e+17, 1.313156379801695e+17, 1.313156379903258e+17, 1.313156380007945e+17, 1.313156380114195e+17, 1.313156380215758e+17, 1.313156380322007e+17, 1.31315638042357e+17, 1.313156380531383e+17, 1.313156380639195e+17, 1.313156380742319e+17, 1.313156380843882e+17, 1.313156380951695e+17, 1.313156381056383e+17, 1.31315638116107e+17, 1.313156381264195e+17, 1.31315638136732e+17, 1.313156381473571e+17, 1.313156381576695e+17, 1.313156381679821e+17, 1.31315638177982e+17, 1.313156381893883e+17, 1.313156382000132e+17, 1.313156382103258e+17, 1.31315638220482e+17, 1.313156382309507e+17, 1.313156382415758e+17, 1.313156382522007e+17, 1.31315638262982e+17, 1.313156382740758e+17, 1.313156382843882e+17, 1.313156382943884e+17, 1.31315638304857e+17, 1.313156383153257e+17, 1.313156383264195e+17, 1.31315638337982e+17, 1.313156383490758e+17, 1.31315638359232e+17, 1.313156383695444e+17, 1.313156383895444e+17, 1.313156384007945e+17, 1.313156384112632e+17, 1.313156384214195e+17, 1.313156384320444e+17, 1.313156384422008e+17, 1.313156384525133e+17, 1.313156384626696e+17, 1.313156384732945e+17, 1.313156384840758e+17, 1.313156384943882e+17, 1.313156385056381e+17, 1.313156385157944e+17, 1.31315638526107e+17, 1.313156385365756e+17, 1.313156385472008e+17, 1.313156385576695e+17, 1.31315638569232e+17, 1.313156385795444e+17, 1.313156385900132e+17, 1.313156386007945e+17, 1.31315638611732e+17, 1.31315638622982e+17, 1.313156386331382e+17, 1.31315638643607e+17, 1.313156386539195e+17, 1.313156386640756e+17, 1.313156386745445e+17, 1.313156386862633e+17, 1.313156386970445e+17, 1.313156387075133e+17, 1.313156387193882e+17, 1.313156387300133e+17, 1.31315638740482e+17, 1.313156387511069e+17, 1.313156387612632e+17, 1.31315638771732e+17, 1.313156387820444e+17, 1.313156387936069e+17, 1.313156388043882e+17, 1.313156388143884e+17, 1.313156388245445e+17, 1.31315638834857e+17, 1.313156388454821e+17, 1.313156388562633e+17, 1.313156388681382e+17, 1.313156388782945e+17, 1.313156388890757e+17, 1.313156388997007e+17, 1.313156389097007e+17, 1.313156389197007e+17, 1.313156389303258e+17, 1.313156389409508e+17, 1.313156389509508e+17, 1.31315638961732e+17, 1.313156389723571e+17, 1.313156389826696e+17, 1.313156389928257e+17, 1.313156390039195e+17, 1.313156390140756e+17, 1.313156390243882e+17, 1.313156390347007e+17, 1.31315639045482e+17, 1.313156390568883e+17, 1.313156390670445e+17, 1.313156390773569e+17, 1.313156390878258e+17, 1.313156390995444e+17, 1.31315639109857e+17, 1.313156391201695e+17, 1.313156391306382e+17, 1.313156391414195e+17, 1.313156391522008e+17, 1.31315639162982e+17, 1.313156391731383e+17, 1.313156391843884e+17, 1.313156391950132e+17, 1.313156392059507e+17, 1.31315639216732e+17, 1.313156392273569e+17, 1.313156392379821e+17, 1.313156392487633e+17, 1.313156392589194e+17, 1.31315639269232e+17, 1.313156392793883e+17, 1.313156392897007e+17, 1.313156393000133e+17, 1.313156393111069e+17, 1.31315639321732e+17, 1.313156393322008e+17, 1.313156393426694e+17, 1.313156393534508e+17, 1.313156393645444e+17, 1.31315639374857e+17, 1.31315639385482e+17, 1.31315639396107e+17, 1.313156394064195e+17, 1.313156394172008e+17, 1.313156394275133e+17, 1.313156394387633e+17, 1.313156394489196e+17, 1.313156394597007e+17, 1.313156394703258e+17, 1.313156394812632e+17, 1.31315639491732e+17, 1.313156395022008e+17, 1.313156395126696e+17, 1.313156395228257e+17, 1.313156395328257e+17, 1.313156395428257e+17, 1.313156395628257e+17, 1.313156395747008e+17, 1.313156395856383e+17, 1.313156395962633e+17, 1.313156396065757e+17, 1.313156396165757e+17, 1.31315639626732e+17, 1.313156396368882e+17, 1.313156396473571e+17, 1.313156396576695e+17, 1.313156396681382e+17, 1.313156396790757e+17, 1.313156396897007e+17, 1.313156397006382e+17, 1.313156397107945e+17, 1.313156397209508e+17, 1.313156397317321e+17, 1.313156397428257e+17, 1.313156397531383e+17, 1.313156397634508e+17, 1.313156397739195e+17, 1.31315639784857e+17, 1.31315639795482e+17, 1.313156398065757e+17, 1.313156398172008e+17, 1.313156398273571e+17, 1.313156398375133e+17, 1.313156398476695e+17, 1.313156398589196e+17, 1.31315639869232e+17, 1.313156398793883e+17, 1.313156398903258e+17, 1.313156399014195e+17, 1.313156399115758e+17, 1.313156399225133e+17, 1.313156399328259e+17, 1.313156399431383e+17, 1.313156399534508e+17, 1.313156399642319e+17, 1.313156399745445e+17, 1.313156399850132e+17, 1.313156399959507e+17, 1.31315640006107e+17, 1.313156400162633e+17, 1.313156400262632e+17, 1.313156400368882e+17, 1.313156400472008e+17, 1.313156400578257e+17, 1.313156400682945e+17, 1.313156400795444e+17, 1.31315640089857e+17, 1.313156401003258e+17, 1.313156401112632e+17, 1.313156401222007e+17, 1.313156401325133e+17, 1.31315640142982e+17, 1.313156401531382e+17, 1.313156401637633e+17, 1.313156401740758e+17, 1.313156401842319e+17, 1.313156401943882e+17, 1.313156402057946e+17, 1.31315640216107e+17, 1.313156402265757e+17, 1.313156402382945e+17, 1.313156402484507e+17, 1.313156402589194e+17, 1.313156402690757e+17, 1.31315640279232e+17, 1.313156402895444e+17, 1.313156403007944e+17, 1.313156403115757e+17, 1.313156403218883e+17, 1.31315640332357e+17, 1.313156403437632e+17, 1.313156403539195e+17, 1.313156403640758e+17, 1.313156403742319e+17, 1.313156403843882e+17, 1.313156403947008e+17, 1.313156404050132e+17, 1.313156404153257e+17, 1.31315640426107e+17, 1.313156404368882e+17, 1.313156404478257e+17, 1.31315640457982e+17, 1.313156404682944e+17, 1.313156404789196e+17, 1.313156404895444e+17, 1.313156405001695e+17, 1.313156405103258e+17, 1.313156405206382e+17, 1.313156405309507e+17, 1.313156405409508e+17, 1.313156405515757e+17, 1.313156405620444e+17, 1.31315640572357e+17, 1.313156405828257e+17, 1.313156405939195e+17, 1.313156406042321e+17, 1.313156406143882e+17, 1.313156406245444e+17, 1.31315640634857e+17, 1.313156406451695e+17, 1.313156406556383e+17, 1.313156406659507e+17, 1.313156406764196e+17, 1.31315640686732e+17, 1.313156406968882e+17, 1.313156407078257e+17, 1.31315640719232e+17, 1.313156407297007e+17, 1.31315640739857e+17, 1.313156407503256e+17, 1.313156407614195e+17, 1.31315640772357e+17, 1.31315640782982e+17, 1.313156407934508e+17, 1.313156408037632e+17, 1.313156408140756e+17, 1.313156408245445e+17, 1.31315640834857e+17, 1.31315640845482e+17, 1.313156408564195e+17, 1.313156408672008e+17, 1.313156408773569e+17, 1.313156408889194e+17, 1.31315640899232e+17, 1.313156409095444e+17, 1.313156409200133e+17, 1.313156409317321e+17, 1.31315640942982e+17, 1.313156409531383e+17, 1.313156409647007e+17, 1.313156409753258e+17, 1.313156409859507e+17, 1.313156409964195e+17, 1.313156410065757e+17, 1.313156410168883e+17, 1.313156410275133e+17, 1.313156410381382e+17, 1.313156410489196e+17, 1.313156410620444e+17, 1.313156410726696e+17, 1.31315641083607e+17, 1.313156410937633e+17, 1.313156411040758e+17, 1.313156411147007e+17, 1.31315641124857e+17, 1.313156411351695e+17, 1.313156411457944e+17, 1.313156411570445e+17, 1.313156411679821e+17, 1.313156411782945e+17, 1.313156411884507e+17, 1.31315641198607e+17, 1.313156412097007e+17, 1.313156412201695e+17, 1.313156412306383e+17, 1.31315641241732e+17, 1.313156412518883e+17, 1.31315641262357e+17, 1.313156412725133e+17, 1.313156412826696e+17, 1.313156412928257e+17, 1.313156413028257e+17, 1.31315641312982e+17, 1.313156413231383e+17, 1.313156413336069e+17, 1.313156413439195e+17, 1.313156413543884e+17, 1.313156413650132e+17, 1.313156413764195e+17, 1.313156413868883e+17, 1.313156413970445e+17, 1.313156414075132e+17, 1.313156414178258e+17, 1.313156414287633e+17, 1.313156414395444e+17, 1.313156414497007e+17, 1.313156414600133e+17, 1.313156414701695e+17, 1.313156414806382e+17, 1.313156414909507e+17, 1.313156415022007e+17, 1.31315641512357e+17, 1.313156415226696e+17, 1.313156415334508e+17, 1.313156415445445e+17, 1.313156415553257e+17, 1.313156415665757e+17, 1.31315641576732e+17, 1.313156415870446e+17, 1.313156415976695e+17, 1.313156416078258e+17, 1.313156416182944e+17, 1.31315641628607e+17, 1.313156416387633e+17, 1.313156416495444e+17, 1.31315641659857e+17, 1.313156416700133e+17, 1.313156416806383e+17, 1.313156416918883e+17, 1.313156417026696e+17, 1.313156417132945e+17, 1.313156417236069e+17, 1.313156417340758e+17, 1.313156417442319e+17, 1.313156417547008e+17, 1.313156417653257e+17, 1.313156417765757e+17, 1.313156417870445e+17, 1.313156417976695e+17, 1.313156418084507e+17, 1.31315641818607e+17, 1.313156418293883e+17, 1.313156418400132e+17, 1.313156418509508e+17, 1.313156418620444e+17, 1.313156418720445e+17, 1.31315641882357e+17, 1.313156418925132e+17, 1.313156419028257e+17, 1.313156419137632e+17, 1.313156419248571e+17, 1.313156419350132e+17, 1.313156419459507e+17, 1.313156419570446e+17, 1.313156419672008e+17, 1.31315641977982e+17, 1.31315641989232e+17, 1.313156419995446e+17, 1.31315642009857e+17, 1.313156420204819e+17, 1.313156420311071e+17, 1.313156420425132e+17, 1.313156420528257e+17, 1.313156420631382e+17, 1.313156420734508e+17, 1.31315642083607e+17, 1.313156420947008e+17, 1.31315642106107e+17, 1.313156421164195e+17, 1.313156421273571e+17, 1.313156421375133e+17, 1.313156421476695e+17, 1.313156421584507e+17, 1.31315642169232e+17, 1.313156421804819e+17, 1.313156421911071e+17, 1.313156422014195e+17, 1.313156422126694e+17, 1.31315642222982e+17, 1.313156422334508e+17, 1.31315642243607e+17, 1.313156422539195e+17, 1.313156422642319e+17, 1.313156422742321e+17, 1.313156422847008e+17, 1.313156422951694e+17, 1.31315642305482e+17, 1.313156423157944e+17, 1.313156423264196e+17, 1.313156423373571e+17, 1.313156423478258e+17, 1.313156423584507e+17, 1.313156423690757e+17, 1.31315642379857e+17, 1.313156423901696e+17, 1.31315642400482e+17, 1.313156424107945e+17, 1.313156424209507e+17, 1.313156424314195e+17, 1.313156424425133e+17, 1.313156424528257e+17, 1.313156424631383e+17, 1.313156424734508e+17, 1.313156424934508e+17, 1.313156425037633e+17, 1.313156425142321e+17, 1.313156425342321e+17, 1.313156425445445e+17, 1.313156425547007e+17, 1.313156425650132e+17, 1.313156425764195e+17, 1.313156425872008e+17, 1.313156425984507e+17, 1.313156426090757e+17, 1.313156426193883e+17, 1.313156426293883e+17, 1.313156426406383e+17, 1.313156426514195e+17, 1.313156426628257e+17, 1.31315642672982e+17, 1.313156426847007e+17, 1.31315642694857e+17, 1.313156427050132e+17, 1.313156427151695e+17, 1.313156427257944e+17, 1.31315642736107e+17, 1.313156427462633e+17, 1.313156427565757e+17, 1.313156427670445e+17, 1.313156427775132e+17, 1.31315642787982e+17, 1.313156427981382e+17, 1.31315642808607e+17, 1.313156428193883e+17, 1.313156428301696e+17, 1.313156428406382e+17, 1.313156428514195e+17, 1.313156428618883e+17, 1.31315642872357e+17, 1.313156428828257e+17, 1.313156428936069e+17, 1.313156429037632e+17, 1.313156429139195e+17, 1.313156429251694e+17, 1.313156429353257e+17, 1.313156429457944e+17, 1.313156429564196e+17, 1.313156429673571e+17, 1.313156429778258e+17, 1.313156429881382e+17, 1.31315642999232e+17, 1.313156430106383e+17, 1.31315643021732e+17, 1.31315643032357e+17, 1.313156430426696e+17, 1.313156430531383e+17, 1.313156430634508e+17, 1.313156430737633e+17, 1.313156430842319e+17, 1.313156430943882e+17, 1.313156431047008e+17, 1.313156431150132e+17, 1.313156431257946e+17, 1.313156431370445e+17, 1.313156431473571e+17, 1.313156431576695e+17, 1.313156431684508e+17, 1.31315643178607e+17, 1.313156431889194e+17, 1.313156431995446e+17, 1.313156432103258e+17, 1.313156432204819e+17, 1.313156432311071e+17, 1.313156432414195e+17, 1.313156432515758e+17, 1.313156432618883e+17, 1.313156432731382e+17, 1.313156432839195e+17, 1.313156432940758e+17, 1.313156433050132e+17, 1.313156433150132e+17, 1.313156433256383e+17, 1.313156433370445e+17, 1.313156433475132e+17, 1.313156433576695e+17, 1.313156433678258e+17, 1.313156433779821e+17, 1.313156433884508e+17, 1.313156433987633e+17, 1.313156434097007e+17, 1.313156434203256e+17, 1.313156434307945e+17, 1.31315643441732e+17, 1.313156434518883e+17, 1.31315643462357e+17, 1.313156434726694e+17, 1.31315643482982e+17, 1.313156434937632e+17, 1.313156435042319e+17, 1.313156435147008e+17, 1.313156435265757e+17, 1.313156435372008e+17, 1.313156435481384e+17, 1.313156435582944e+17, 1.313156435684508e+17, 1.313156435790758e+17, 1.313156435893883e+17, 1.313156435997007e+17, 1.313156436100133e+17, 1.313156436203258e+17, 1.313156436306382e+17, 1.313156436418883e+17, 1.313156436522007e+17, 1.313156436626694e+17, 1.313156436731382e+17, 1.313156436832945e+17, 1.313156436934508e+17, 1.31315643703607e+17, 1.313156437137632e+17, 1.313156437240756e+17, 1.313156437351695e+17, 1.31315643745482e+17, 1.31315643756107e+17, 1.313156437675133e+17, 1.313156437781382e+17, 1.313156437893883e+17, 1.313156437997007e+17, 1.313156438101695e+17, 1.31315643820482e+17, 1.313156438312634e+17, 1.313156438415758e+17, 1.31315643851732e+17, 1.31315643862982e+17, 1.31315643873607e+17, 1.313156438837632e+17, 1.313156438940756e+17, 1.313156439051694e+17, 1.313156439157946e+17, 1.313156439264195e+17, 1.31315643936732e+17, 1.313156439468883e+17, 1.313156439573569e+17, 1.313156439679821e+17, 1.313156439784508e+17, 1.313156439890757e+17, 1.31315643999857e+17, 1.31315644010482e+17, 1.313156440212632e+17, 1.313156440315757e+17, 1.313156440425133e+17, 1.313156440526694e+17, 1.313156440632945e+17, 1.313156440734508e+17, 1.313156440836069e+17, 1.313156440942321e+17, 1.31315644104857e+17, 1.31315644115482e+17, 1.31315644126107e+17, 1.313156441370445e+17, 1.313156441475132e+17, 1.313156441576695e+17, 1.313156441687633e+17, 1.313156441790757e+17, 1.31315644189857e+17, 1.313156442000133e+17, 1.313156442114195e+17, 1.313156442228257e+17, 1.313156442340758e+17, 1.313156442442321e+17, 1.313156442545445e+17, 1.31315644264857e+17, 1.313156442750132e+17, 1.31315644285482e+17, 1.313156442956383e+17, 1.31315644306107e+17, 1.313156443165757e+17, 1.313156443268883e+17, 1.313156443376695e+17, 1.313156443481382e+17, 1.313156443582944e+17, 1.313156443684507e+17, 1.313156443793883e+17, 1.313156443903258e+17, 1.313156444007945e+17, 1.313156444111069e+17, 1.313156444212632e+17, 1.313156444318883e+17, 1.313156444422007e+17, 1.31315644452357e+17, 1.313156444625133e+17, 1.31315644472982e+17, 1.313156444832945e+17, 1.31315644493607e+17, 1.313156445042321e+17, 1.313156445147008e+17, 1.313156445264195e+17, 1.313156445372008e+17, 1.313156445478257e+17, 1.313156445589196e+17, 1.31315644569232e+17, 1.313156445795444e+17, 1.313156445897007e+17, 1.313156446000133e+17, 1.313156446101696e+17, 1.31315644620482e+17, 1.313156446309508e+17, 1.313156446415758e+17, 1.313156446522007e+17, 1.31315644662982e+17, 1.313156446736069e+17, 1.313156446942319e+17, 1.313156447043882e+17, 1.313156447145445e+17, 1.313156447247007e+17, 1.313156447351695e+17, 1.313156447457944e+17, 1.313156447564196e+17, 1.313156447665756e+17, 1.313156447778258e+17, 1.313156447879821e+17, 1.313156447990757e+17, 1.31315644809232e+17, 1.31315644819857e+17, 1.313156448312634e+17, 1.31315644841732e+17, 1.31315644852357e+17, 1.313156448625132e+17, 1.31315644873607e+17, 1.313156448840758e+17, 1.313156448943884e+17, 1.313156449047008e+17, 1.313156449151695e+17, 1.313156449257944e+17, 1.313156449364195e+17, 1.31315644946732e+17, 1.313156449570445e+17, 1.313156449673571e+17, 1.31315644977982e+17, 1.313156449881382e+17, 1.313156449984507e+17, 1.313156450087633e+17, 1.313156450189196e+17, 1.313156450293883e+17, 1.313156450397007e+17, 1.313156450500133e+17, 1.313156450601696e+17, 1.313156450706382e+17, 1.313156450807945e+17, 1.313156450915757e+17, 1.313156451026696e+17, 1.313156451134508e+17, 1.313156451237632e+17, 1.313156451340758e+17, 1.313156451443882e+17, 1.313156451550132e+17, 1.313156451656383e+17, 1.313156451759507e+17, 1.313156451872008e+17, 1.313156451984507e+17, 1.31315645208607e+17, 1.313156452189196e+17, 1.313156452290757e+17, 1.313156452393883e+17, 1.313156452497007e+17, 1.31315645259857e+17, 1.313156452703258e+17, 1.313156452806382e+17, 1.313156452907945e+17, 1.313156453015758e+17, 1.313156453118883e+17, 1.313156453225133e+17, 1.313156453337633e+17, 1.313156453440758e+17, 1.313156453547007e+17, 1.313156453650132e+17, 1.313156453756383e+17, 1.313156453856383e+17, 1.313156453962633e+17, 1.313156454068882e+17, 1.313156454176695e+17, 1.31315645427982e+17, 1.313156454381382e+17, 1.313156454481382e+17, 1.313156454587633e+17, 1.313156454690758e+17, 1.313156454797007e+17, 1.313156454909508e+17, 1.313156455012634e+17, 1.313156455114195e+17, 1.313156455215757e+17, 1.313156455325133e+17, 1.313156455426696e+17, 1.313156455532945e+17, 1.313156455637633e+17, 1.313156455745445e+17, 1.313156455847008e+17, 1.313156455950132e+17, 1.313156456050132e+17, 1.31315645615482e+17, 1.313156456267319e+17, 1.313156456373571e+17, 1.313156456489196e+17, 1.313156456601695e+17, 1.313156456703258e+17, 1.31315645680482e+17, 1.313156456911069e+17, 1.313156457015757e+17, 1.31315645711732e+17, 1.313156457226694e+17, 1.313156457331382e+17, 1.313156457432945e+17, 1.313156457540758e+17, 1.313156457642321e+17, 1.313156457750132e+17, 1.313156457859507e+17, 1.313156457962633e+17, 1.313156458065757e+17, 1.313156458176695e+17, 1.31315645827982e+17, 1.313156458381382e+17, 1.313156458482945e+17, 1.313156458584508e+17, 1.31315645869232e+17, 1.313156458795444e+17, 1.313156458897007e+17, 1.313156459000133e+17, 1.313156459109508e+17, 1.313156459212632e+17, 1.313156459312632e+17, 1.313156459418883e+17, 1.313156459522007e+17, 1.313156459626694e+17, 1.313156459731382e+17, 1.313156459832945e+17, 1.313156459934508e+17, 1.313156460037633e+17, 1.313156460142319e+17, 1.313156460245445e+17, 1.313156460350132e+17, 1.313156460450132e+17, 1.313156460564195e+17, 1.313156460672008e+17, 1.313156460776695e+17, 1.313156460884507e+17, 1.31315646099232e+17, 1.313156461093883e+17, 1.313156461197007e+17, 1.313156461300133e+17, 1.313156461401695e+17, 1.313156461504819e+17, 1.313156461606382e+17, 1.313156461714195e+17, 1.313156461815758e+17, 1.31315646192357e+17, 1.31315646202982e+17, 1.313156462140758e+17, 1.313156462242321e+17, 1.313156462345445e+17, 1.313156462445445e+17, 1.313156462545445e+17, 1.313156462647007e+17, 1.313156462750132e+17, 1.313156462851695e+17, 1.313156462956381e+17, 1.313156463057944e+17, 1.313156463164195e+17, 1.313156463265757e+17, 1.313156463365757e+17, 1.313156463470445e+17, 1.313156463572008e+17, 1.313156463681384e+17, 1.31315646378607e+17, 1.313156463887633e+17, 1.31315646399232e+17, 1.31315646409857e+17, 1.313156464203258e+17, 1.313156464304819e+17, 1.313156464411071e+17, 1.313156464512632e+17, 1.313156464614195e+17, 1.31315646471732e+17, 1.313156464822007e+17, 1.313156464926696e+17, 1.313156465039195e+17, 1.313156465140758e+17, 1.313156465243884e+17, 1.313156465347008e+17, 1.31315646544857e+17, 1.31315646555482e+17, 1.313156465668883e+17, 1.313156465775132e+17, 1.313156465878257e+17, 1.31315646597982e+17, 1.313156466084507e+17, 1.313156466187633e+17, 1.313156466293883e+17, 1.313156466400133e+17, 1.313156466503258e+17, 1.31315646660482e+17, 1.313156466707945e+17, 1.313156466814194e+17, 1.313156466914195e+17, 1.313156467020444e+17, 1.313156467131383e+17, 1.313156467237632e+17, 1.313156467340758e+17, 1.313156467442321e+17, 1.313156467545445e+17, 1.313156467647007e+17, 1.313156467751695e+17, 1.313156467853257e+17, 1.313156467957946e+17, 1.313156468078257e+17, 1.313156468178258e+17, 1.313156468279821e+17, 1.313156468389196e+17, 1.313156468490757e+17, 1.31315646859232e+17, 1.313156468700133e+17, 1.313156468801695e+17, 1.313156468903258e+17, 1.313156469015758e+17, 1.313156469122007e+17, 1.313156469228257e+17, 1.31315646932982e+17, 1.31315646943607e+17, 1.313156469540758e+17, 1.313156469642321e+17, 1.313156469747007e+17, 1.313156469857944e+17, 1.313156469959507e+17, 1.313156470065757e+17, 1.31315647016732e+17, 1.31315647026732e+17, 1.313156470370445e+17, 1.313156470482945e+17, 1.31315647058607e+17, 1.313156470689194e+17, 1.313156470793882e+17, 1.313156470900133e+17, 1.313156471001696e+17, 1.313156471103258e+17, 1.31315647120482e+17, 1.313156471307945e+17, 1.313156471412632e+17, 1.313156471515757e+17, 1.313156471625132e+17, 1.313156471732945e+17, 1.31315647183607e+17, 1.313156471940756e+17, 1.313156472042321e+17, 1.313156472147008e+17, 1.313156472251694e+17, 1.313156472357944e+17, 1.313156472465757e+17, 1.313156472567319e+17, 1.313156472670445e+17, 1.313156472773569e+17, 1.313156472879821e+17, 1.313156472987633e+17, 1.313156473095444e+17, 1.313156473203258e+17, 1.313156473311071e+17, 1.31315647341732e+17, 1.313156473523571e+17, 1.313156473626696e+17, 1.313156473726694e+17, 1.313156473832946e+17, 1.313156473937632e+17, 1.313156474042321e+17, 1.313156474143884e+17, 1.31315647424857e+17, 1.31315647436107e+17, 1.313156474464196e+17, 1.31315647456732e+17, 1.313156474672008e+17, 1.31315647477982e+17, 1.313156474882945e+17, 1.313156474984507e+17, 1.31315647508607e+17, 1.313156475187633e+17, 1.313156475290757e+17, 1.313156475398569e+17, 1.313156475503258e+17, 1.313156475609508e+17, 1.313156475717321e+17, 1.313156475820445e+17, 1.313156475926694e+17, 1.313156476028257e+17, 1.313156476132945e+17, 1.313156476237632e+17, 1.313156476340758e+17, 1.313156476447008e+17, 1.313156476550132e+17, 1.313156476653258e+17, 1.313156476756383e+17, 1.31315647686107e+17, 1.313156476972006e+17, 1.313156477078258e+17, 1.313156477178257e+17, 1.313156477284508e+17, 1.313156477389194e+17, 1.313156477495446e+17, 1.313156477597007e+17, 1.313156477701695e+17, 1.313156477812632e+17, 1.313156477915758e+17, 1.31315647802357e+17, 1.313156478128257e+17, 1.313156478234508e+17, 1.313156478337632e+17, 1.313156478450132e+17, 1.313156478553258e+17, 1.31315647865482e+17, 1.313156478756383e+17, 1.313156478859507e+17, 1.313156478968882e+17, 1.313156479078258e+17, 1.313156479182944e+17, 1.313156479284507e+17, 1.313156479387633e+17, 1.313156479489196e+17, 1.313156479590757e+17, 1.313156479695444e+17, 1.313156479797007e+17, 1.313156479900132e+17, 1.313156480007945e+17, 1.313156480111071e+17, 1.313156480217321e+17, 1.31315648031732e+17, 1.313156480425133e+17, 1.31315648052982e+17, 1.313156480634508e+17, 1.31315648073607e+17, 1.313156480842319e+17, 1.313156480943882e+17, 1.313156481047008e+17, 1.313156481151694e+17, 1.313156481259507e+17, 1.31315648136107e+17, 1.313156481464196e+17, 1.313156481568882e+17, 1.313156481681382e+17, 1.313156481781382e+17, 1.313156481890757e+17, 1.313156481997007e+17, 1.313156482104819e+17, 1.313156482214195e+17, 1.313156482322008e+17, 1.313156482423571e+17, 1.313156482526696e+17, 1.313156482631383e+17, 1.313156482740758e+17, 1.313156482842321e+17, 1.313156482947008e+17, 1.313156483051695e+17, 1.313156483151695e+17, 1.31315648326107e+17, 1.313156483375132e+17, 1.313156483475132e+17, 1.313156483578258e+17, 1.313156483687633e+17, 1.31315648379857e+17, 1.313156483901695e+17, 1.313156484009508e+17, 1.313156484112632e+17, 1.313156484214195e+17, 1.313156484318883e+17, 1.313156484422008e+17, 1.313156484525133e+17, 1.313156484628259e+17, 1.313156484732945e+17, 1.313156484843882e+17, 1.313156484947007e+17, 1.313156485050132e+17, 1.313156485162633e+17, 1.313156485264195e+17, 1.31315648536732e+17, 1.313156485470445e+17, 1.313156485573569e+17, 1.313156485676695e+17, 1.31315648578607e+17, 1.313156485887633e+17, 1.313156485995444e+17, 1.313156486100133e+17, 1.313156486203258e+17, 1.313156486312632e+17, 1.313156486414195e+17, 1.313156486515757e+17, 1.313156486625133e+17, 1.313156486728257e+17, 1.313156486828257e+17, 1.313156486931383e+17, 1.31315648703607e+17, 1.313156487142319e+17, 1.313156487243882e+17, 1.313156487347008e+17, 1.313156487450132e+17, 1.31315648756732e+17, 1.313156487673571e+17, 1.313156487776695e+17, 1.313156487881382e+17, 1.313156487987633e+17, 1.313156488090758e+17, 1.313156488197007e+17, 1.31315648830482e+17, 1.313156488412632e+17, 1.31315648851732e+17, 1.31315648861732e+17, 1.313156488720444e+17, 1.313156488828257e+17, 1.31315648892982e+17, 1.313156489031382e+17, 1.313156489134508e+17, 1.31315648923607e+17, 1.313156489340756e+17, 1.313156489450132e+17, 1.31315648955482e+17, 1.313156489659508e+17, 1.313156489765757e+17, 1.313156489868882e+17, 1.313156489972008e+17, 1.31315649007982e+17, 1.313156490182945e+17, 1.313156490284508e+17, 1.313156490390757e+17, 1.313156490501695e+17, 1.313156490604819e+17, 1.313156490711069e+17, 1.313156490812632e+17, 1.313156490922008e+17, 1.31315649102982e+17, 1.313156491132945e+17, 1.313156491236069e+17, 1.313156491337632e+17, 1.313156491442319e+17, 1.313156491547008e+17, 1.313156491650132e+17, 1.31315649175482e+17, 1.313156491864196e+17, 1.313156491975132e+17, 1.313156492076695e+17, 1.313156492182944e+17, 1.31315649229232e+17, 1.313156492395444e+17, 1.313156492493882e+17, 1.313156492603258e+17, 1.31315649270482e+17, 1.31315649280482e+17, 1.313156492903258e+17, 1.313156493003258e+17, 1.313156493103258e+17, 1.31315649321732e+17, 1.31315649332357e+17, 1.313156493432945e+17, 1.31315649353607e+17, 1.313156493639195e+17, 1.313156493739195e+17, 1.313156493836069e+17, 1.313156493931383e+17, 1.31315649402357e+17, 1.313156494120445e+17, 1.313156494218883e+17, 1.313156494307945e+17, 1.313156494409508e+17, 1.313156494500133e+17, 1.313156494595444e+17, 1.313156494687633e+17, 1.313156494779821e+17, 1.31315649487982e+17, 1.313156494981382e+17, 1.31315649509232e+17, 1.313156495181382e+17, 1.313156495275132e+17, 1.313156495368883e+17, 1.313156495468883e+17, 1.313156495562633e+17, 1.313156495657944e+17, 1.313156495751695e+17, 1.313156495847007e+17, 1.31315649593607e+17, 1.313156496039195e+17, 1.313156496132945e+17, 1.31315649622357e+17, 1.313156496318883e+17, 1.313156496409508e+17, 1.313156496501695e+17, 1.313156496593882e+17, 1.313156496695444e+17, 1.313156496789194e+17, 1.313156496882945e+17, 1.313156496978258e+17, 1.31315649707982e+17, 1.313156497195444e+17, 1.313156497300133e+17, 1.313156497412632e+17, 1.31315649751732e+17, 1.313156497620444e+17, 1.313156497726696e+17, 1.313156497839195e+17, 1.313156497942319e+17, 1.313156498051695e+17, 1.313156498157946e+17, 1.313156498265757e+17, 1.313156498372008e+17, 1.313156498484507e+17, 1.313156498590757e+17, 1.31315649870482e+17, 1.313156498815757e+17, 1.313156498922007e+17, 1.313156499036069e+17, 1.313156499153258e+17, 1.313156499262633e+17, 1.313156499370445e+17, 1.313156499476695e+17, 1.313156499582944e+17, 1.313156499690757e+17, 1.31315649980482e+17, 1.313156499911069e+17, 1.313156500022008e+17, 1.313156500134508e+17, 1.31315650024857e+17, 1.313156500356383e+17, 1.313156500464195e+17, 1.313156500570445e+17, 1.313156500676695e+17, 1.313156500778257e+17, 1.313156500881382e+17, 1.313156500982945e+17, 1.313156501086071e+17, 1.313156501190757e+17, 1.313156501306383e+17, 1.313156501414195e+17, 1.313156501515757e+17, 1.31315650161732e+17, 1.313156501718883e+17, 1.31315650182357e+17, 1.313156501926696e+17, 1.31315650203607e+17, 1.313156502139195e+17, 1.313156502245445e+17, 1.313156502347007e+17, 1.313156502456383e+17, 1.313156502564195e+17, 1.313156502668882e+17, 1.31315650277982e+17, 1.313156502893882e+17, 1.313156503012632e+17, 1.313156503132946e+17, 1.313156503256383e+17, 1.313156503384507e+17, 1.313156503512632e+17, 1.313156503639195e+17, 1.313156503762632e+17, 1.313156503882945e+17, 1.313156504004819e+17, 1.313156504125133e+17, 1.313156504245445e+17, 1.313156504368883e+17, 1.31315650449232e+17, 1.313156504618883e+17, 1.313156504739195e+17, 1.31315650486107e+17, 1.313156504982945e+17, 1.313156505106382e+17, 1.313156505228257e+17, 1.31315650534857e+17, 1.313156505473571e+17, 1.313156505593883e+17, 1.313156505715758e+17, 1.31315650583607e+17, 1.313156505962632e+17, 1.313156506089196e+17, 1.313156506211069e+17, 1.313156506332945e+17, 1.313156506453257e+17, 1.313156506573571e+17, 1.313156506693883e+17, 1.313156506814195e+17, 1.313156506934508e+17, 1.31315650705482e+17, 1.313156507184508e+17, 1.313156507312634e+17, 1.31315650743607e+17, 1.313156507559507e+17, 1.31315650767982e+17, 1.313156507801695e+17, 1.31315650792357e+17, 1.313156508045445e+17, 1.313156508168883e+17, 1.313156508290757e+17, 1.313156508412634e+17, 1.313156508532945e+17, 1.31315650865482e+17, 1.313156508778258e+17, 1.313156508903258e+17, 1.313156509025133e+17, 1.313156509145445e+17, 1.313156509268883e+17, 1.313156509389196e+17, 1.313156509514195e+17, 1.313156509639195e+17, 1.31315650976107e+17, 1.313156509881382e+17, 1.313156510007945e+17, 1.313156510129819e+17, 1.313156510251695e+17, 1.313156510375133e+17, 1.313156510495446e+17, 1.313156510620444e+17, 1.313156510742319e+17, 1.31315651086732e+17, 1.313156510990757e+17, 1.313156511114195e+17, 1.31315651123607e+17, 1.313156511356383e+17, 1.313156511481382e+17, 1.31315651160482e+17, 1.313156511726694e+17, 1.31315651184857e+17, 1.313156511972008e+17, 1.313156512093883e+17, 1.31315651221732e+17, 1.313156512343884e+17, 1.313156512465757e+17, 1.313156512587633e+17, 1.313156512711069e+17, 1.313156512834508e+17, 1.31315651295482e+17, 1.313156513078258e+17, 1.31315651320482e+17, 1.31315651332982e+17, 1.313156513451694e+17, 1.313156513575132e+17, 1.31315651369857e+17, 1.313156513820445e+17, 1.313156513940758e+17, 1.313156514064196e+17, 1.313156514189196e+17, 1.313156514309507e+17, 1.313156514432945e+17, 1.313156514559507e+17, 1.31315651467982e+17, 1.313156514803258e+17, 1.31315651492357e+17, 1.313156515043882e+17, 1.31315651516732e+17, 1.313156515287633e+17, 1.313156515409508e+17, 1.31315651552982e+17, 1.313156515650132e+17, 1.313156515772008e+17, 1.313156515900132e+17, 1.313156516020445e+17, 1.313156516147008e+17, 1.31315651626732e+17, 1.313156516387633e+17, 1.313156516507945e+17, 1.313156516628257e+17, 1.313156516748571e+17, 1.313156516872008e+17, 1.313156516995444e+17, 1.313156517117321e+17, 1.313156517242319e+17, 1.313156517362633e+17, 1.313156517487633e+17, 1.313156517607944e+17, 1.313156517732945e+17, 1.313156517853258e+17, 1.313156517973571e+17, 1.313156518095446e+17, 1.313156518218883e+17, 1.313156518340758e+17, 1.31315651846107e+17, 1.313156518582945e+17, 1.313156518703258e+17, 1.313156518826694e+17, 1.31315651894857e+17, 1.313156519068883e+17, 1.313156519193882e+17, 1.313156519320444e+17, 1.31315651944857e+17, 1.313156519568883e+17, 1.313156519693883e+17, 1.313156519815758e+17, 1.31315651993607e+17, 1.313156520059508e+17, 1.313156520179821e+17, 1.313156520301696e+17, 1.31315652042357e+17, 1.313156520543884e+17, 1.313156520665757e+17, 1.313156520790757e+17, 1.313156520912632e+17, 1.313156521034508e+17, 1.31315652115482e+17, 1.313156521275132e+17, 1.313156521397007e+17, 1.313156521518883e+17, 1.313156521639195e+17, 1.31315652176107e+17, 1.313156521884507e+17, 1.31315652200482e+17, 1.313156522125133e+17, 1.31315652224857e+17, 1.313156522368882e+17, 1.31315652249232e+17, 1.313156522615758e+17, 1.313156522739195e+17, 1.313156522859507e+17, 1.313156522979821e+17, 1.313156523103258e+17, 1.313156523223571e+17, 1.313156523347008e+17, 1.31315652346732e+17, 1.313156523590757e+17, 1.313156523714195e+17, 1.313156523837633e+17, 1.313156523957946e+17, 1.313156524079821e+17, 1.313156524201695e+17, 1.31315652432357e+17, 1.313156524445445e+17, 1.313156524565757e+17, 1.31315652468607e+17, 1.313156524807945e+17, 1.313156524931383e+17, 1.313156525057946e+17, 1.313156525179821e+17, 1.31315652530482e+17, 1.313156525425133e+17, 1.313156525545445e+17, 1.31315652566732e+17, 1.313156525789196e+17, 1.313156525914195e+17, 1.31315652603607e+17, 1.313156526157946e+17, 1.313156526281382e+17, 1.313156526403258e+17, 1.31315652652357e+17, 1.313156526647008e+17, 1.31315652676732e+17, 1.313156526887633e+17, 1.313156527009508e+17, 1.313156527134508e+17, 1.313156527256383e+17, 1.313156527378258e+17, 1.313156527503258e+17, 1.31315652762357e+17, 1.313156527743882e+17, 1.313156527865757e+17, 1.313156527987633e+17, 1.313156528109508e+17, 1.31315652822982e+17, 1.313156528353257e+17, 1.313156528475132e+17, 1.313156528597007e+17, 1.31315652871732e+17, 1.313156528837632e+17, 1.313156528962632e+17, 1.31315652908607e+17, 1.313156529207945e+17, 1.313156529328257e+17, 1.31315652945482e+17, 1.313156529575132e+17, 1.313156529697007e+17, 1.31315652981732e+17, 1.313156529937632e+17, 1.31315653006107e+17, 1.313156530187633e+17, 1.313156530307945e+17, 1.313156530426694e+17, 1.313156530547007e+17, 1.31315653066732e+17, 1.313156530787633e+17, 1.313156530907945e+17, 1.313156531028257e+17},
			             {1.313156411147007e+17, 1.31315641124857e+17, 1.313156411351695e+17, 1.313156411457944e+17},
			             {1.313156376500132e+17, 1.313156376615758e+17, 1.313156376722007e+17, 1.31315637682357e+17, 1.313156376926694e+17, 1.313156377034508e+17, 1.31315637713607e+17, 1.313156377237632e+17, 1.313156377347007e+17, 1.313156377451695e+17, 1.313156377557944e+17, 1.31315637766107e+17, 1.313156377776695e+17, 1.313156377881382e+17, 1.313156377984507e+17, 1.313156378093883e+17, 1.313156378211071e+17, 1.31315637831732e+17, 1.313156382415758e+17, 1.313156382843882e+17, 1.31315638304857e+17, 1.313156383153257e+17, 1.31315638337982e+17, 1.313156383490758e+17, 1.313156383695444e+17, 1.313156384112632e+17, 1.313156384214195e+17, 1.313156384320444e+17, 1.313156384422008e+17, 1.313156384626696e+17, 1.313156384732945e+17, 1.313156385056381e+17, 1.313156385157944e+17, 1.31315638526107e+17, 1.313156385365756e+17, 1.313156385472008e+17, 1.313156385795444e+17, 1.313156385900132e+17, 1.31315638611732e+17, 1.31315638622982e+17, 1.313156386539195e+17, 1.313156386640756e+17, 1.313156386862633e+17, 1.313156386970445e+17, 1.313156387193882e+17, 1.313156387300133e+17, 1.31315639269232e+17, 1.313156392793883e+17, 1.313156392897007e+17, 1.313156393000133e+17, 1.31315639626732e+17, 1.313156396368882e+17, 1.313156396473571e+17, 1.313156396576695e+17, 1.313156396681382e+17, 1.313156396790757e+17, 1.313156396897007e+17, 1.313156397006382e+17, 1.313156397107945e+17, 1.313156397317321e+17, 1.313156397428257e+17, 1.313156397531383e+17, 1.313156397634508e+17, 1.313156397739195e+17, 1.31315639784857e+17, 1.31315639795482e+17, 1.313156398065757e+17, 1.313156398172008e+17, 1.313156398273571e+17, 1.313156398375133e+17, 1.313156398476695e+17, 1.313156398589196e+17, 1.31315639869232e+17, 1.313156398793883e+17, 1.313156398903258e+17, 1.313156399014195e+17, 1.313156399115758e+17, 1.313156399225133e+17, 1.313156399328259e+17, 1.313156399431383e+17, 1.313156399534508e+17, 1.313156399642319e+17, 1.313156399745445e+17, 1.313156399850132e+17, 1.313156399959507e+17, 1.313156400162633e+17, 1.313156400262632e+17, 1.313156400682945e+17, 1.313156403539195e+17, 1.313156403640758e+17, 1.313156403742319e+17, 1.313156403843882e+17, 1.313156403947008e+17, 1.313156404050132e+17, 1.313156404153257e+17, 1.31315640426107e+17, 1.313156404368882e+17, 1.313156404478257e+17, 1.31315640457982e+17, 1.313156404682944e+17, 1.313156404789196e+17, 1.313156404895444e+17, 1.313156405001695e+17, 1.313156405103258e+17, 1.313156405206382e+17, 1.313156405309507e+17, 1.313156405409508e+17, 1.313156405515757e+17, 1.313156405620444e+17, 1.31315640572357e+17, 1.313156405828257e+17, 1.313156405939195e+17, 1.313156406042321e+17, 1.313156406143882e+17, 1.313156406245444e+17, 1.31315640634857e+17, 1.313156406451695e+17, 1.313156406556383e+17, 1.313156406659507e+17, 1.313156406764196e+17, 1.31315640686732e+17, 1.313156406968882e+17, 1.313156407078257e+17, 1.31315640719232e+17, 1.313156407297007e+17, 1.31315640739857e+17, 1.313156407503256e+17, 1.313156407614195e+17, 1.31315640772357e+17, 1.31315640782982e+17, 1.313156407934508e+17, 1.313156408037632e+17, 1.313156408140756e+17, 1.313156408245445e+17, 1.31315640834857e+17, 1.31315640845482e+17, 1.313156408564195e+17, 1.313156408672008e+17, 1.313156408773569e+17, 1.313156408889194e+17, 1.31315640899232e+17, 1.313156409095444e+17, 1.313156409200133e+17, 1.313156409317321e+17, 1.31315640942982e+17, 1.313156409531383e+17, 1.313156409647007e+17, 1.313156409753258e+17, 1.313156409859507e+17, 1.313156409964195e+17, 1.313156410065757e+17, 1.313156410168883e+17, 1.313156410275133e+17, 1.313156410381382e+17, 1.313156410489196e+17, 1.313156410620444e+17, 1.313156410726696e+17, 1.31315641083607e+17, 1.313156410937633e+17, 1.313156411040758e+17, 1.313156411147007e+17, 1.31315641124857e+17, 1.313156411351695e+17, 1.313156411457944e+17, 1.313156411570445e+17, 1.313156411679821e+17, 1.313156411782945e+17, 1.313156411884507e+17, 1.31315641198607e+17, 1.313156412097007e+17, 1.313156412201695e+17, 1.313156412306383e+17, 1.31315641241732e+17, 1.313156412518883e+17, 1.31315641262357e+17, 1.313156412725133e+17, 1.313156412826696e+17, 1.313156412928257e+17, 1.313156413028257e+17, 1.31315641312982e+17, 1.313156413231383e+17, 1.313156413336069e+17, 1.313156413439195e+17, 1.313156413543884e+17, 1.313156413650132e+17, 1.313156413764195e+17, 1.313156413868883e+17, 1.313156413970445e+17, 1.313156414075132e+17, 1.313156414178258e+17, 1.313156414287633e+17, 1.313156414395444e+17, 1.313156414497007e+17, 1.313156414600133e+17, 1.313156414701695e+17, 1.313156414806382e+17, 1.313156414909507e+17, 1.313156415022007e+17, 1.31315641512357e+17, 1.313156415226696e+17, 1.313156415334508e+17, 1.313156415445445e+17, 1.313156415553257e+17, 1.313156415665757e+17, 1.31315641576732e+17, 1.313156415870446e+17, 1.313156415976695e+17, 1.313156416078258e+17, 1.313156416182944e+17, 1.313156416387633e+17, 1.313156416495444e+17, 1.31315641659857e+17, 1.313156416700133e+17, 1.313156416806383e+17, 1.313156416918883e+17, 1.313156417026696e+17, 1.313156417132945e+17, 1.313156417236069e+17, 1.313156417340758e+17, 1.313156417442319e+17, 1.313156417547008e+17, 1.313156417653257e+17, 1.313156417765757e+17, 1.313156417870445e+17, 1.313156417976695e+17, 1.313156418084507e+17, 1.31315641818607e+17, 1.313156418293883e+17, 1.313156418400132e+17, 1.313156418509508e+17, 1.313156418620444e+17, 1.313156418720445e+17, 1.31315641882357e+17, 1.313156418925132e+17, 1.313156419028257e+17, 1.313156419137632e+17, 1.313156419248571e+17, 1.313156419350132e+17, 1.313156419459507e+17, 1.313156419570446e+17, 1.313156419672008e+17, 1.31315641977982e+17, 1.31315641989232e+17, 1.313156419995446e+17, 1.31315642009857e+17, 1.313156420204819e+17, 1.313156420311071e+17, 1.313156420425132e+17, 1.313156420528257e+17, 1.313156420631382e+17, 1.313156420734508e+17, 1.31315642083607e+17, 1.313156420947008e+17, 1.31315642106107e+17, 1.313156421273571e+17, 1.313156421375133e+17, 1.313156421476695e+17, 1.313156421584507e+17, 1.31315642169232e+17, 1.313156421804819e+17, 1.313156421911071e+17, 1.313156422014195e+17, 1.313156422126694e+17, 1.31315642222982e+17, 1.313156422334508e+17, 1.31315642243607e+17, 1.313156422539195e+17, 1.313156422642319e+17, 1.313156422742321e+17, 1.313156422847008e+17, 1.313156422951694e+17, 1.31315642305482e+17, 1.313156423157944e+17, 1.313156423264196e+17, 1.313156423373571e+17, 1.313156423478258e+17, 1.313156423584507e+17, 1.313156423690757e+17, 1.31315642379857e+17, 1.313156423901696e+17, 1.31315642400482e+17, 1.313156424107945e+17, 1.313156424209507e+17, 1.313156424314195e+17, 1.313156424425133e+17, 1.313156424528257e+17, 1.313156424631383e+17, 1.313156424734508e+17, 1.313156424934508e+17, 1.313156425037633e+17, 1.313156425142321e+17, 1.313156425342321e+17, 1.313156425445445e+17, 1.313156425547007e+17, 1.313156425650132e+17, 1.313156425764195e+17, 1.313156425872008e+17, 1.313156425984507e+17, 1.313156426090757e+17, 1.313156426193883e+17, 1.313156426293883e+17, 1.313156426406383e+17, 1.313156426514195e+17, 1.313156426628257e+17, 1.31315642672982e+17, 1.313156426847007e+17, 1.31315642694857e+17, 1.313156427151695e+17, 1.313156427565757e+17, 1.31315642808607e+17, 1.313156428514195e+17, 1.31315643032357e+17, 1.313156430426696e+17, 1.313156430531383e+17, 1.313156430634508e+17, 1.313156430737633e+17, 1.313156430842319e+17, 1.313156430943882e+17, 1.313156431047008e+17, 1.313156431150132e+17, 1.313156431257946e+17, 1.313156431370445e+17, 1.313156431473571e+17, 1.313156431576695e+17, 1.313156431684508e+17, 1.31315643178607e+17, 1.313156431889194e+17, 1.313156431995446e+17, 1.313156432103258e+17, 1.313156432204819e+17, 1.313156432311071e+17, 1.313156432414195e+17, 1.313156432515758e+17, 1.313156432618883e+17, 1.313156432731382e+17, 1.313156432839195e+17, 1.313156432940758e+17, 1.313156433050132e+17, 1.313156433150132e+17, 1.313156433256383e+17, 1.313156433370445e+17, 1.313156433475132e+17, 1.313156433576695e+17, 1.313156433678258e+17, 1.313156433779821e+17, 1.313156433884508e+17, 1.313156433987633e+17, 1.313156434097007e+17, 1.313156434203256e+17, 1.313156434307945e+17, 1.31315643441732e+17, 1.313156434518883e+17, 1.31315643462357e+17, 1.313156434726694e+17, 1.31315643482982e+17, 1.313156434937632e+17, 1.313156435042319e+17, 1.313156435147008e+17, 1.313156435265757e+17, 1.313156435372008e+17, 1.313156435582944e+17, 1.313156435684508e+17, 1.313156435790758e+17, 1.313156435893883e+17, 1.313156435997007e+17, 1.313156436100133e+17, 1.313156436203258e+17, 1.313156436306382e+17, 1.313156436418883e+17, 1.313156436522007e+17, 1.313156436832945e+17, 1.31315643703607e+17, 1.313156437137632e+17, 1.313156437240756e+17, 1.313156437351695e+17, 1.31315643745482e+17, 1.313156437675133e+17, 1.313156437893883e+17, 1.313156437997007e+17, 1.313156438101695e+17, 1.31315643820482e+17, 1.313156438312634e+17, 1.313156438415758e+17, 1.31315643851732e+17, 1.31315643862982e+17, 1.31315643873607e+17, 1.313156438837632e+17, 1.313156438940756e+17, 1.313156439051694e+17, 1.313156439157946e+17, 1.313156439264195e+17, 1.31315643936732e+17, 1.313156439468883e+17, 1.313156439573569e+17, 1.313156439679821e+17, 1.313156439784508e+17, 1.313156439890757e+17, 1.31315643999857e+17, 1.31315644010482e+17, 1.313156440212632e+17, 1.313156440315757e+17, 1.313156440425133e+17, 1.313156440526694e+17, 1.313156440632945e+17, 1.313156440734508e+17, 1.313156440942321e+17, 1.31315644104857e+17, 1.31315644115482e+17, 1.31315644126107e+17, 1.313156441370445e+17, 1.313156441475132e+17, 1.313156441576695e+17, 1.313156441687633e+17, 1.313156441790757e+17, 1.31315644189857e+17, 1.313156442000133e+17, 1.313156442114195e+17, 1.313156442228257e+17, 1.313156442340758e+17, 1.313156442442321e+17, 1.313156442545445e+17, 1.31315644264857e+17, 1.313156442750132e+17, 1.31315644285482e+17, 1.313156442956383e+17, 1.31315644306107e+17, 1.313156443165757e+17, 1.313156443268883e+17, 1.313156443376695e+17, 1.313156443481382e+17, 1.313156443582944e+17, 1.313156443684507e+17, 1.313156443793883e+17, 1.313156443903258e+17, 1.313156444007945e+17, 1.313156444111069e+17, 1.313156444212632e+17, 1.313156444318883e+17, 1.313156444422007e+17, 1.31315644452357e+17, 1.313156444625133e+17, 1.31315644472982e+17, 1.313156444832945e+17, 1.31315644493607e+17, 1.313156445042321e+17, 1.313156445147008e+17, 1.313156445264195e+17, 1.313156445372008e+17, 1.313156445478257e+17, 1.313156445589196e+17, 1.31315644569232e+17, 1.313156445795444e+17, 1.313156445897007e+17, 1.313156446000133e+17, 1.313156446101696e+17, 1.31315644620482e+17, 1.313156446309508e+17, 1.313156446415758e+17, 1.313156446522007e+17, 1.31315644662982e+17, 1.313156446736069e+17, 1.313156446942319e+17, 1.313156447043882e+17, 1.313156447145445e+17, 1.313156447247007e+17, 1.313156447351695e+17, 1.313156447457944e+17, 1.313156447564196e+17, 1.313156447665756e+17, 1.313156447778258e+17, 1.313156447879821e+17, 1.313156447990757e+17, 1.31315644809232e+17, 1.31315644819857e+17, 1.313156448312634e+17, 1.31315644841732e+17, 1.31315644852357e+17, 1.313156448625132e+17, 1.31315644873607e+17, 1.313156448840758e+17, 1.313156448943884e+17, 1.313156449047008e+17, 1.313156449151695e+17, 1.313156449257944e+17, 1.313156449364195e+17, 1.31315644946732e+17, 1.313156449570445e+17, 1.313156449673571e+17, 1.31315644977982e+17, 1.313156449881382e+17, 1.313156449984507e+17, 1.313156450087633e+17, 1.313156450189196e+17, 1.313156450397007e+17, 1.313156450500133e+17, 1.313156450601696e+17, 1.313156452703258e+17, 1.313156452806382e+17, 1.313156453547007e+17, 1.313156453650132e+17, 1.313156453756383e+17, 1.313156453856383e+17, 1.313156453962633e+17, 1.313156454068882e+17, 1.313156454176695e+17, 1.31315645427982e+17, 1.313156454381382e+17, 1.313156454481382e+17, 1.313156454587633e+17, 1.313156454690758e+17, 1.313156454797007e+17, 1.313156454909508e+17, 1.313156455012634e+17, 1.313156455114195e+17, 1.313156455215757e+17, 1.313156455325133e+17, 1.313156455426696e+17, 1.313156455532945e+17, 1.313156455637633e+17, 1.313156455745445e+17, 1.313156455847008e+17, 1.313156455950132e+17, 1.313156456050132e+17, 1.31315645615482e+17, 1.313156456267319e+17, 1.313156456373571e+17, 1.313156456489196e+17, 1.313156456601695e+17, 1.313156456703258e+17, 1.31315645680482e+17, 1.313156456911069e+17, 1.313156457015757e+17, 1.31315645711732e+17, 1.313156457226694e+17, 1.313156457331382e+17, 1.313156457432945e+17, 1.313156457540758e+17, 1.313156457642321e+17, 1.313156457750132e+17, 1.313156457859507e+17, 1.313156457962633e+17, 1.313156458065757e+17, 1.313156458176695e+17, 1.31315645827982e+17, 1.313156458381382e+17, 1.313156458482945e+17, 1.313156458584508e+17, 1.31315645869232e+17, 1.313156458795444e+17, 1.313156458897007e+17, 1.313156459000133e+17, 1.313156463470445e+17, 1.313156463572008e+17, 1.313156463681384e+17, 1.31315646399232e+17, 1.31315646409857e+17, 1.313156464304819e+17, 1.313156464411071e+17, 1.313156464614195e+17, 1.31315646471732e+17, 1.313156464822007e+17, 1.313156464926696e+17, 1.313156465039195e+17, 1.313156465140758e+17, 1.313156465347008e+17, 1.31315646544857e+17, 1.31315646555482e+17, 1.313156465668883e+17, 1.313156465775132e+17, 1.313156465878257e+17, 1.31315646597982e+17, 1.313156466084507e+17, 1.313156466187633e+17, 1.313156466293883e+17, 1.313156466400133e+17, 1.313156466503258e+17, 1.31315646660482e+17, 1.313156466707945e+17, 1.313156466814194e+17, 1.313156466914195e+17, 1.313156467131383e+17, 1.313156467442321e+17, 1.313156467545445e+17, 1.313156467647007e+17, 1.313156467751695e+17, 1.313156467853257e+17, 1.313156467957946e+17, 1.313156468279821e+17, 1.313156468389196e+17, 1.313156468490757e+17, 1.31315646859232e+17, 1.313156468801695e+17, 1.313156468903258e+17, 1.313156469015758e+17, 1.313156469122007e+17, 1.31315646932982e+17, 1.31315646943607e+17, 1.313156469857944e+17, 1.313156469959507e+17, 1.31315647016732e+17, 1.31315647026732e+17, 1.313156470482945e+17, 1.31315647058607e+17, 1.313156470793882e+17, 1.313156470900133e+17, 1.313156471515757e+17, 1.313156471625132e+17, 1.313156471940756e+17, 1.313156472042321e+17, 1.313156472357944e+17, 1.313156472465757e+17, 1.313156472773569e+17, 1.313156472879821e+17, 1.313156473203258e+17, 1.313156473311071e+17, 1.313156474672008e+17, 1.31315647477982e+17, 1.313156475290757e+17, 1.313156475398569e+17, 1.313156475926694e+17, 1.313156476028257e+17, 1.313156476447008e+17, 1.313156476550132e+17, 1.313156477078258e+17, 1.313156477178257e+17, 1.313156477701695e+17, 1.313156477812632e+17, 1.313156478234508e+17, 1.313156478337632e+17, 1.313156483578258e+17, 1.313156483687633e+17, 1.313156484628259e+17, 1.313156484732945e+17, 1.313156485676695e+17, 1.31315648578607e+17, 1.313156486625133e+17, 1.313156486728257e+17, 1.313156487243882e+17, 1.313156487347008e+17, 1.313156488197007e+17, 1.31315648830482e+17, 1.313156489134508e+17, 1.31315648923607e+17, 1.31315649007982e+17, 1.313156490182945e+17, 1.313156490812632e+17, 1.313156490922008e+17, 1.313156491650132e+17, 1.31315649175482e+17, 1.313156492493882e+17, 1.313156492603258e+17, 1.313156493432945e+17, 1.31315649353607e+17, 1.313156493836069e+17, 1.313156493931383e+17, 1.313156494687633e+17, 1.313156494779821e+17, 1.313156495468883e+17, 1.313156495562633e+17, 1.31315649622357e+17, 1.313156496318883e+17, 1.313156496882945e+17, 1.313156496978258e+17, 1.313156497620444e+17, 1.313156497726696e+17, 1.313156498372008e+17, 1.313156498484507e+17, 1.313156499153258e+17, 1.313156499262633e+17, 1.313156499911069e+17, 1.313156500022008e+17, 1.313156500356383e+17, 1.313156500464195e+17, 1.313156500778257e+17, 1.313156500881382e+17, 1.313156501306383e+17, 1.313156501414195e+17, 1.313156501718883e+17, 1.31315650182357e+17, 1.313156502139195e+17, 1.313156502245445e+17, 1.313156502668882e+17, 1.31315650277982e+17, 1.313156503132946e+17, 1.313156503256383e+17, 1.313156503639195e+17, 1.313156503762632e+17, 1.313156504125133e+17, 1.313156504245445e+17, 1.313156504618883e+17, 1.313156504739195e+17, 1.313156504982945e+17, 1.313156505106382e+17, 1.313156505473571e+17, 1.313156505593883e+17, 1.313156506089196e+17, 1.313156506211069e+17, 1.313156506573571e+17, 1.313156506693883e+17, 1.31315650705482e+17, 1.313156507184508e+17, 1.313156507559507e+17, 1.31315650767982e+17, 1.313156508045445e+17, 1.313156508168883e+17, 1.313156508532945e+17, 1.31315650865482e+17, 1.313156508778258e+17, 1.313156509025133e+17, 1.313156509145445e+17, 1.313156509389196e+17, 1.313156509514195e+17, 1.313156509639195e+17, 1.31315650976107e+17, 1.313156510251695e+17, 1.313156510375133e+17, 1.313156510742319e+17, 1.31315651086732e+17, 1.313156510990757e+17, 1.313156511114195e+17, 1.31315651123607e+17, 1.313156511356383e+17, 1.313156511481382e+17, 1.31315651160482e+17, 1.313156511726694e+17, 1.31315651184857e+17, 1.313156511972008e+17, 1.313156512093883e+17, 1.31315651221732e+17, 1.313156512343884e+17, 1.313156512465757e+17, 1.313156512587633e+17, 1.313156512711069e+17, 1.313156512834508e+17, 1.31315651295482e+17, 1.313156513078258e+17, 1.31315651320482e+17, 1.31315651332982e+17, 1.313156513451694e+17, 1.313156513575132e+17, 1.31315651369857e+17, 1.313156513820445e+17, 1.313156513940758e+17, 1.313156514064196e+17, 1.313156514189196e+17, 1.313156514309507e+17, 1.313156514432945e+17, 1.313156514559507e+17, 1.31315651467982e+17, 1.313156514803258e+17, 1.31315651492357e+17, 1.313156515043882e+17, 1.31315651516732e+17, 1.313156515287633e+17, 1.313156515409508e+17, 1.31315651552982e+17, 1.313156515650132e+17, 1.313156515772008e+17, 1.313156515900132e+17, 1.313156516020445e+17, 1.313156516147008e+17, 1.31315651626732e+17, 1.313156516387633e+17, 1.313156516507945e+17, 1.313156516628257e+17, 1.313156516748571e+17, 1.313156516872008e+17, 1.313156516995444e+17, 1.313156517117321e+17, 1.313156517242319e+17, 1.313156517362633e+17, 1.313156517487633e+17, 1.313156517607944e+17, 1.313156517732945e+17, 1.313156517853258e+17, 1.313156517973571e+17, 1.313156518095446e+17, 1.313156518218883e+17, 1.313156518340758e+17, 1.31315651846107e+17, 1.313156518582945e+17, 1.313156518703258e+17, 1.313156518826694e+17, 1.31315651894857e+17, 1.313156519068883e+17, 1.313156519193882e+17, 1.313156519320444e+17, 1.31315651944857e+17, 1.313156519568883e+17, 1.313156519693883e+17, 1.313156519815758e+17, 1.31315651993607e+17, 1.313156520059508e+17, 1.313156520179821e+17, 1.313156520301696e+17, 1.31315652042357e+17, 1.313156520543884e+17, 1.313156520665757e+17, 1.313156520790757e+17, 1.313156520912632e+17, 1.313156521034508e+17, 1.31315652115482e+17, 1.313156521275132e+17, 1.313156521397007e+17, 1.313156521518883e+17, 1.313156521639195e+17, 1.31315652176107e+17, 1.313156521884507e+17, 1.31315652200482e+17, 1.313156522125133e+17, 1.31315652224857e+17, 1.313156522368882e+17, 1.31315652249232e+17, 1.313156522615758e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
