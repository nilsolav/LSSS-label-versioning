netcdf mask {
	:date_created = "20200811T114915";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200811T114915";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 21;
			channels = 6;
			categories = 126;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  21.2, 20.7, 19.9, 24.3, 19.2, 17.3, 18.8, 18.6, 27.2, 27.1, 35.5, 25.9, 28.9, 33.6, 28.8,  2.4, 63.1,  3.9, 64.3, 20.2, 38.6;
			max_depth =  34.6, 34.5, 24.9, 31.2, 25.9, 31.7, 24.7, 34.7, 35.8, 34.7, 46.6, 38.8, 43.8, 37.8, 43.6,  2.8, 66.3,  4.1, 67.7, 22.5, 45.2;
			start_time = 131376817067200768, 131376811774388224, 131376811962669440, 131376812029857024, 131376812074388224, 131376812235169536, 131376812638607104, 131376812893294464, 131376818492669568, 131376819050169472, 131376825916732032, 131376827864700800, 131376828991419520, 131376829317981952, 131376829617200768, 131376828167981952, 131376827970794496, 131376832800794496, 131376825672513280, 131376821250638336, 131376832738294400;
			end_time = 131376817115638272, 131376811839544448, 131376811987044480, 131376812040169600, 131376812092825728, 131376812289232000, 131376812651419520, 131376812930325760, 131376818552669568, 131376819063607040, 131376825996107008, 131376827911888256, 131376829102044544, 131376829332513280, 131376829838138240, 131376828167981952, 131376828010638208, 131376832800794496, 131376825712982016, 131376821254857088, 131376832770638208;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "6009", "6009", "6009", "6009", "6009", "6009", "5027", "5027", "5027", "5027", "5027", "5027", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "6009", "6009", "6009", "6009", "6009", "6009", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "6009", "6009", "6009", "6009", "6009", "6009", "1", "1", "1", "1", "1", "1", "6009", "6009", "6009", "6009", "6009", "6009", "0", "0", "0", "0", "0", "0", "1", "1", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63;
			mask_times = {1.313768170672008e+17, 1.313768171156383e+17},
			             {1.313768117743882e+17, 1.313768118395444e+17},
			             {1.313768119626694e+17, 1.313768119870445e+17},
			             {1.31376812029857e+17, 1.313768120401696e+17},
			             {1.313768120743882e+17, 1.313768120928257e+17},
			             {1.313768122351695e+17, 1.31376812289232e+17},
			             {1.313768126386071e+17, 1.313768126514195e+17},
			             {1.313768128932945e+17, 1.313768129303258e+17},
			             {1.313768184926696e+17, 1.313768185526696e+17},
			             {1.313768190501695e+17, 1.31376819063607e+17},
			             {1.31376825916732e+17, 1.31376825996107e+17},
			             {1.313768278647008e+17, 1.313768279118883e+17},
			             {1.313768289914195e+17, 1.313768291020445e+17},
			             {1.31376829317982e+17, 1.313768293325133e+17},
			             {1.313768296172008e+17, 1.313768296265757e+17, 1.313768296364195e+17, 1.313768296407945e+17, 1.31376829650482e+17, 1.313768296597009e+17, 1.313768296640758e+17, 1.313768296734508e+17, 1.31376829683607e+17, 1.313768296878258e+17, 1.313768297025133e+17, 1.313768297126696e+17, 1.313768297226694e+17, 1.313768297273571e+17, 1.313768297370445e+17, 1.31376829746732e+17, 1.313768297515758e+17, 1.313768297614195e+17, 1.313768297656383e+17, 1.313768297712632e+17, 1.313768297840756e+17, 1.313768298381382e+17},
			             {1.31376828167982e+17},
			             {1.313768279707945e+17, 1.313768280106382e+17},
			             {1.313768328007945e+17},
			             {1.313768256725133e+17, 1.31376825712982e+17},
			             {1.313768212506383e+17, 1.313768212548571e+17},
			             {1.313768327382944e+17, 1.313768327706382e+17};
			mask_depths = {{21.2, 34.6}, {21.2, 34.6}}, {{20.7, 34.5}, {20.7, 34.5}}, {{19.9, 24.9}, {19.9, 24.9}}, {{24.3, 31.2}, {24.3, 31.2}}, {{19.2, 25.9}, {19.2, 25.9}}, {{17.3, 31.7}, {17.3, 31.7}}, {{18.8, 24.7}, {18.8, 24.7}}, {{18.6, 34.7}, {18.6, 34.7}}, {{27.2, 35.8}, {27.2, 35.8}}, {{27.1, 34.7}, {27.1, 34.7}}, {{35.5, 46.6}, {35.5, 46.6}}, {{25.9, 38.8}, {25.9, 38.8}}, {{28.9, 43.8}, {28.9, 43.8}}, {{33.6, 37.8}, {33.6, 37.8}}, {{37.8, 40.6, 40.8}, {36.3, 37.7, 40.5}, {36.0, 36.2}, {35.6, 35.9, 40.7, 40.9}, {35.1, 35.5, 41.0, 41.3}, {34.5, 35.0, 41.4, 41.5}, {33.9, 34.4}, {33.3, 33.8, 41.7, 42.2}, {32.8, 33.2, 42.3, 42.4}, {32.2, 32.7, 42.5, 43.3}, {43.4, 43.5}, {43.6}, {31.8, 31.9}, {31.6, 31.7}, {31.1, 31.5}, {30.7, 31.0}, {30.4, 30.6}, {30.0, 30.3}, {29.6, 29.9}, {28.8, 28.9, 29.5}, {29.0}, {29.0, 43.6}}, {{2.4, 2.4, 2.8, 2.8}}, {{63.1, 66.3}, {63.1, 66.3}}, {{3.9, 3.9, 4.1, 4.1}}, {{64.3, 67.7}, {64.3, 67.7}}, {{20.2, 22.5}, {20.2, 22.5}}, {{38.6, 45.2}, {38.6, 45.2}};
		}
	}
}
