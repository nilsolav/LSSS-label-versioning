netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 43;
			channels = 6;
			categories = 258;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0,  9.6, 63.1, 14.0, 13.9, 61.2, 55.5, 60.3, 62.7, 64.2, 65.3, 64.1, 68.2, 32.7, 31.9, 65.3, 52.3, 53.9, 54.1, 62.8, 52.5, 52.9, 56.9, 54.7, 51.0, 55.3, 57.4, 49.6, 58.5, 55.5, 60.5, 68.6, 68.0, 60.4, 64.8, 61.4, 62.3, 11.2, 10.9,  9.8, 11.6, 61.2, 64.2;
			max_depth =  65.6, 76.7, 64.4, 26.9, 23.9, 65.0, 61.4, 62.3, 65.7, 65.8, 66.7, 65.8, 69.2, 35.8, 34.0, 72.3, 61.7, 66.7, 58.6, 68.4, 60.6, 54.0, 60.3, 57.8, 62.4, 64.7, 62.2, 57.2, 64.1, 61.8, 67.8, 69.7, 69.7, 63.1, 67.3, 63.9, 64.9, 31.3, 31.8, 31.9, 34.4, 63.2, 65.7;
			start_time = 128874387948804480, 128874389460835712, 128874388596773248, 128874400233209600, 128874400761334528, 128874398341334528, 128874401549303168, 128874402789303296, 128874402801334528, 128874395088804480, 128874391672867072, 128874392076773248, 128874393788804608, 128874397881334528, 128874395220835840, 128874406385240704, 128874408653209600, 128874409037272064, 128874409289303296, 128874409405240704, 128874409773209472, 128874409837272064, 128874410841334400, 128874410957271936, 128874412153209472, 128874412605240832, 128874414613209472, 128874415501334528, 128874416701334400, 128874417641334528, 128874420469303296, 128874416169303296, 128874421789303296, 128874428217271936, 128874422545240832, 128874427081334528, 128874430521334528, 128874425541334528, 128874425693209472, 128874430621334528, 128874432065240704, 128874423169303168, 128874423381334400;
			end_time = 128874389460835712, 128874435034569600, 128874388620835840, 128874400465240832, 128874401045240704, 128874398365240832, 128874401573209472, 128874402805240704, 128874402829303296, 128874395112866944, 128874391696773248, 128874392092867072, 128874393808804480, 128874397901334400, 128874395236773248, 128874406449303296, 128874408741334528, 128874409221334528, 128874409353209472, 128874409449303168, 128874409833209472, 128874409853209472, 128874410861334528, 128874410989303296, 128874412261334528, 128874412665240832, 128874414661334400, 128874415585240704, 128874416733209472, 128874417693209472, 128874420521334400, 128874416197272064, 128874421833209472, 128874428253209472, 128874422581334528, 128874427117272064, 128874430549303168, 128874425677271936, 128874426753209472, 128874430841334528, 128874432413209472, 128874423193209472, 128874423417271936;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43;
			region_name = "Layer1","Layer2","Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21","Layer22","Layer23","Layer24","Layer25","Layer26","Layer27","Layer28","Layer29","Layer30","Layer31","Layer32","Layer33","Layer34","Layer35","Layer36","Layer37","Layer38","Layer39","Layer40","Layer41";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63;
			mask_times = {1.288743879488045e+17, 1.288743879528669e+17, 1.288743879567732e+17, 1.288743879608357e+17, 1.288743879648983e+17, 1.288743879688045e+17, 1.288743879728671e+17, 1.288743879767732e+17, 1.288743879808357e+17, 1.288743879848983e+17, 1.288743879888045e+17, 1.288743879928669e+17, 1.288743879967732e+17, 1.288743880008357e+17, 1.288743880048983e+17, 1.288743880088045e+17, 1.288743880128671e+17, 1.288743880167732e+17, 1.288743880208357e+17, 1.288743880248983e+17, 1.288743880288045e+17, 1.288743880328671e+17, 1.288743880367731e+17, 1.288743880408357e+17, 1.288743880448983e+17, 1.288743880488045e+17, 1.288743880528671e+17, 1.288743880567732e+17, 1.288743880608357e+17, 1.288743880648983e+17, 1.288743880688045e+17, 1.288743880728671e+17, 1.288743880767732e+17, 1.288743880808357e+17, 1.288743880848983e+17, 1.288743880888045e+17, 1.288743880928671e+17, 1.288743880967732e+17, 1.288743881008358e+17, 1.288743881048983e+17, 1.288743881088045e+17, 1.288743881128671e+17, 1.288743881167732e+17, 1.288743881208357e+17, 1.288743881248982e+17, 1.288743881288045e+17, 1.288743881328671e+17, 1.288743881367732e+17, 1.288743881408358e+17, 1.288743881448982e+17, 1.288743881488045e+17, 1.288743881528669e+17, 1.288743881567732e+17, 1.288743881608358e+17, 1.288743881648982e+17, 1.288743881688045e+17, 1.288743881728669e+17, 1.288743881767732e+17, 1.288743881808357e+17, 1.288743881848983e+17, 1.288743881888046e+17, 1.288743881928669e+17, 1.288743881967732e+17, 1.288743882008357e+17, 1.288743882048982e+17, 1.288743882088045e+17, 1.288743882128669e+17, 1.288743882167732e+17, 1.288743882208357e+17, 1.288743882248983e+17, 1.288743882288045e+17, 1.288743882328671e+17, 1.288743882367732e+17, 1.288743882408357e+17, 1.288743882448983e+17, 1.288743882488045e+17, 1.288743882528669e+17, 1.288743882567732e+17, 1.288743882608357e+17, 1.288743882648983e+17, 1.288743882688045e+17, 1.288743882728671e+17, 1.288743882767732e+17, 1.288743882808357e+17, 1.288743882848983e+17, 1.288743882888045e+17, 1.288743882928671e+17, 1.288743882967731e+17, 1.288743883008357e+17, 1.288743883048983e+17, 1.288743883088045e+17, 1.288743883128671e+17, 1.288743883167732e+17, 1.288743883208357e+17, 1.288743883248983e+17, 1.288743883288045e+17, 1.288743883328671e+17, 1.288743883367732e+17, 1.288743883408357e+17, 1.288743883448983e+17, 1.288743883488045e+17, 1.288743883528671e+17, 1.288743883567732e+17, 1.288743883608358e+17, 1.288743883648982e+17, 1.288743883688045e+17, 1.288743883728671e+17, 1.288743883767732e+17, 1.288743883808357e+17, 1.288743883848982e+17, 1.288743883888045e+17, 1.288743883928669e+17, 1.288743883967732e+17, 1.288743884008358e+17, 1.288743884048983e+17, 1.288743884088045e+17, 1.288743884128669e+17, 1.288743884167732e+17, 1.288743884208357e+17, 1.288743884248982e+17, 1.288743884288045e+17, 1.288743884328669e+17, 1.288743884367732e+17, 1.288743884408357e+17, 1.288743884448983e+17, 1.288743884488045e+17, 1.288743884528669e+17, 1.288743884567732e+17, 1.288743884608357e+17, 1.288743884648983e+17, 1.288743884688045e+17, 1.288743884728669e+17, 1.288743884767732e+17, 1.288743884808357e+17, 1.288743884848983e+17, 1.288743884888045e+17, 1.288743884928671e+17, 1.288743884967732e+17, 1.288743885008357e+17, 1.288743885048983e+17, 1.288743885088045e+17, 1.288743885128669e+17, 1.288743885167732e+17, 1.288743885208357e+17, 1.288743885248983e+17, 1.288743885288045e+17, 1.288743885328671e+17, 1.288743885367732e+17, 1.288743885408357e+17, 1.288743885448983e+17, 1.288743885488045e+17, 1.288743885528671e+17, 1.288743885567732e+17, 1.288743885608357e+17, 1.288743885648983e+17, 1.288743885688045e+17, 1.288743885728671e+17, 1.288743885767732e+17, 1.288743885808357e+17, 1.288743885848983e+17, 1.288743885888045e+17, 1.288743885928671e+17, 1.288743885967732e+17, 1.288743886008357e+17, 1.288743886048983e+17, 1.288743886088045e+17, 1.288743886128671e+17, 1.288743886167732e+17, 1.288743886208358e+17, 1.288743886248982e+17, 1.288743886288045e+17, 1.288743886328671e+17, 1.288743886367732e+17, 1.288743886408357e+17, 1.288743886448982e+17, 1.288743886488045e+17, 1.288743886528669e+17, 1.288743886567732e+17, 1.288743886608358e+17, 1.288743886648983e+17, 1.288743886688045e+17, 1.288743886728669e+17, 1.288743886767732e+17, 1.288743886808357e+17, 1.288743886848982e+17, 1.288743886888045e+17, 1.288743886928669e+17, 1.288743886967732e+17, 1.288743887008357e+17, 1.288743887048983e+17, 1.288743887088045e+17, 1.288743887128669e+17, 1.288743887167732e+17, 1.288743887208357e+17, 1.288743887248983e+17, 1.288743887288045e+17, 1.288743887328669e+17, 1.288743887367732e+17, 1.288743887408357e+17, 1.288743887448983e+17, 1.288743887488045e+17, 1.288743887528671e+17, 1.288743887567732e+17, 1.288743887608357e+17, 1.288743887648983e+17, 1.288743887688045e+17, 1.288743887728669e+17, 1.288743887767732e+17, 1.288743887808357e+17, 1.288743887848983e+17, 1.288743887888045e+17, 1.288743887928671e+17, 1.288743887967732e+17, 1.288743888008357e+17, 1.288743888048983e+17, 1.288743888088045e+17, 1.288743888128671e+17, 1.288743888167732e+17, 1.288743888208357e+17, 1.288743888248983e+17, 1.288743888288045e+17, 1.288743888328671e+17, 1.288743888367732e+17, 1.288743888408357e+17, 1.288743888448983e+17, 1.288743888488045e+17, 1.288743888528671e+17, 1.288743888567732e+17, 1.288743888608357e+17, 1.288743888648983e+17, 1.288743888688045e+17, 1.288743888728671e+17, 1.288743888767732e+17, 1.288743888808358e+17, 1.288743888848982e+17, 1.288743888888045e+17, 1.288743888928671e+17, 1.288743888967732e+17, 1.288743889008357e+17, 1.288743889048982e+17, 1.288743889088045e+17, 1.288743889128669e+17, 1.288743889167732e+17, 1.288743889208358e+17, 1.288743889248983e+17, 1.288743889288046e+17, 1.288743889328669e+17, 1.288743889367732e+17, 1.288743889408357e+17, 1.288743889448982e+17, 1.288743889488045e+17, 1.288743889528669e+17, 1.288743889567732e+17, 1.288743889608357e+17, 1.288743889648983e+17, 1.288743889688045e+17, 1.288743889728669e+17, 1.288743889767732e+17, 1.288743889808357e+17, 1.288743889848983e+17, 1.288743889888045e+17, 1.288743889928669e+17, 1.288743889967732e+17, 1.288743890008357e+17, 1.288743890048983e+17, 1.288743890088045e+17, 1.288743890128671e+17, 1.288743890167732e+17, 1.288743890208357e+17, 1.288743890248983e+17, 1.288743890288045e+17, 1.288743890328669e+17, 1.288743890367732e+17, 1.288743890408357e+17, 1.288743890448983e+17, 1.288743890488045e+17, 1.288743890528671e+17, 1.288743890567732e+17, 1.288743890608357e+17, 1.288743890648983e+17, 1.288743890688045e+17, 1.288743890728671e+17, 1.288743890767732e+17, 1.288743890808357e+17, 1.288743890848983e+17, 1.288743890888045e+17, 1.288743890928671e+17, 1.288743890967732e+17, 1.288743891008357e+17, 1.288743891048983e+17, 1.288743891088045e+17, 1.288743891128671e+17, 1.288743891167732e+17, 1.288743891208357e+17, 1.288743891248982e+17, 1.288743891288045e+17, 1.288743891328671e+17, 1.288743891367732e+17, 1.288743891408358e+17, 1.288743891448982e+17, 1.288743891488045e+17, 1.288743891528671e+17, 1.288743891567732e+17, 1.288743891608357e+17, 1.288743891648982e+17, 1.288743891688045e+17, 1.288743891728669e+17, 1.288743891767732e+17, 1.288743891808358e+17, 1.288743891848983e+17, 1.288743891888046e+17, 1.288743891928669e+17, 1.288743891967732e+17, 1.288743892008357e+17, 1.288743892048982e+17, 1.288743892088045e+17, 1.288743892128669e+17, 1.288743892167732e+17, 1.288743892208357e+17, 1.288743892248983e+17, 1.288743892288045e+17, 1.288743892328669e+17, 1.288743892367732e+17, 1.288743892408357e+17, 1.288743892448983e+17, 1.288743892488045e+17, 1.288743892528669e+17, 1.288743892567732e+17, 1.288743892608357e+17, 1.288743892648983e+17, 1.288743892688045e+17, 1.288743892728671e+17, 1.288743892767732e+17, 1.288743892808357e+17, 1.288743892848983e+17, 1.288743892888045e+17, 1.288743892928669e+17, 1.288743892967732e+17, 1.288743893008357e+17, 1.288743893048983e+17, 1.288743893088045e+17, 1.288743893128671e+17, 1.288743893167732e+17, 1.288743893208357e+17, 1.288743893248983e+17, 1.288743893288045e+17, 1.288743893328671e+17, 1.288743893367732e+17, 1.288743893408357e+17, 1.288743893448983e+17, 1.288743893488045e+17, 1.288743893528671e+17, 1.288743893567732e+17, 1.288743893608358e+17, 1.288743893648983e+17, 1.288743893688045e+17, 1.288743893728671e+17, 1.288743893767732e+17, 1.288743893808357e+17, 1.288743893848982e+17, 1.288743893888045e+17, 1.288743893928671e+17, 1.288743893967732e+17, 1.288743894008358e+17, 1.288743894048982e+17, 1.288743894088045e+17, 1.288743894128669e+17, 1.288743894167732e+17, 1.288743894208357e+17, 1.288743894248982e+17, 1.288743894288045e+17, 1.288743894328669e+17, 1.288743894367732e+17, 1.288743894408357e+17, 1.288743894448983e+17, 1.288743894488046e+17, 1.288743894528669e+17, 1.288743894567732e+17, 1.288743894608357e+17},
			             {1.288743894608357e+17, 1.288743894648982e+17, 1.288743894688045e+17, 1.288743894728669e+17, 1.288743894767732e+17, 1.288743894808357e+17, 1.288743894848983e+17, 1.288743894888045e+17, 1.288743894928669e+17, 1.288743894967732e+17, 1.288743895008357e+17, 1.288743895048983e+17, 1.288743895088045e+17, 1.288743895128669e+17, 1.288743895167732e+17, 1.288743895208357e+17, 1.288743895248983e+17, 1.288743895288045e+17, 1.288743895328671e+17, 1.288743895367732e+17, 1.288743895408357e+17, 1.288743895448983e+17, 1.288743895488045e+17, 1.288743895528669e+17, 1.288743895567732e+17, 1.288743895608357e+17, 1.288743895648983e+17, 1.288743895688045e+17, 1.288743895728671e+17, 1.288743895767732e+17, 1.288743895808357e+17, 1.288743895848983e+17, 1.288743895888045e+17, 1.288743895928671e+17, 1.288743895967732e+17, 1.288743896008357e+17, 1.288743896048983e+17, 1.288743896088045e+17, 1.288743896128671e+17, 1.288743896167732e+17, 1.288743896208358e+17, 1.288743896248983e+17, 1.288743896288045e+17, 1.288743896328671e+17, 1.288743896367732e+17, 1.288743896408357e+17, 1.288743896448982e+17, 1.288743896488045e+17, 1.288743896528671e+17, 1.288743896567732e+17, 1.288743896608358e+17, 1.288743896648982e+17, 1.288743896688045e+17, 1.288743896728669e+17, 1.288743896767732e+17, 1.288743896808358e+17, 1.288743896848982e+17, 1.288743896888045e+17, 1.288743896928669e+17, 1.288743896967732e+17, 1.288743897008357e+17, 1.288743897048983e+17, 1.288743897088046e+17, 1.288743897128669e+17, 1.288743897167732e+17, 1.288743897208357e+17, 1.288743897248982e+17, 1.288743897288045e+17, 1.288743897328669e+17, 1.288743897367732e+17, 1.288743897408357e+17, 1.288743897448983e+17, 1.288743897488045e+17, 1.288743897528671e+17, 1.288743897567732e+17, 1.288743897608357e+17, 1.288743897648983e+17, 1.288743897688045e+17, 1.288743897728669e+17, 1.288743897767732e+17, 1.288743897808357e+17, 1.288743897848983e+17, 1.288743897888045e+17, 1.288743897928671e+17, 1.288743897967732e+17, 1.288743898008357e+17, 1.288743898048983e+17, 1.288743898088045e+17, 1.288743898128671e+17, 1.288743898167731e+17, 1.288743898208357e+17, 1.288743898248983e+17, 1.288743898288045e+17, 1.288743898328671e+17, 1.288743898367732e+17, 1.288743898408357e+17, 1.288743898448983e+17, 1.288743898488045e+17, 1.288743898528671e+17, 1.288743898567732e+17, 1.288743898608357e+17, 1.288743898648983e+17, 1.288743898688045e+17, 1.288743898728671e+17, 1.288743898767732e+17, 1.288743898808358e+17, 1.288743898848983e+17, 1.288743898888045e+17, 1.288743898928671e+17, 1.288743898967732e+17, 1.288743899008357e+17, 1.288743899048982e+17, 1.288743899088045e+17, 1.288743899128671e+17, 1.288743899167732e+17, 1.288743899208358e+17, 1.288743899248982e+17, 1.288743899288045e+17, 1.288743899328669e+17, 1.288743899367732e+17, 1.288743899408358e+17, 1.288743899448982e+17, 1.288743899488045e+17, 1.288743899528669e+17, 1.288743899567732e+17, 1.288743899608357e+17, 1.288743899648983e+17, 1.288743899688046e+17, 1.288743899728669e+17, 1.288743899767732e+17, 1.288743899808357e+17, 1.288743899848982e+17, 1.288743899888045e+17, 1.288743899928669e+17, 1.288743899967732e+17, 1.288743900008357e+17, 1.288743900048983e+17, 1.288743900088045e+17, 1.288743900128671e+17, 1.288743900167732e+17, 1.288743900208357e+17, 1.288743900248983e+17, 1.288743900288045e+17, 1.288743900328669e+17, 1.288743900367732e+17, 1.288743900408357e+17, 1.288743900448983e+17, 1.288743900488045e+17, 1.288743900528671e+17, 1.288743900567732e+17, 1.288743900608357e+17, 1.288743900648983e+17, 1.288743900688045e+17, 1.288743900728671e+17, 1.288743900767731e+17, 1.288743900808357e+17, 1.288743900848983e+17, 1.288743900888045e+17, 1.288743900928671e+17, 1.288743900967732e+17, 1.288743901008357e+17, 1.288743901048983e+17, 1.288743901088045e+17, 1.288743901128671e+17, 1.288743901167732e+17, 1.288743901208357e+17, 1.288743901248983e+17, 1.288743901288045e+17, 1.288743901328671e+17, 1.288743901367732e+17, 1.288743901408358e+17, 1.288743901448982e+17, 1.288743901488045e+17, 1.288743901528671e+17, 1.288743901567732e+17, 1.288743901608357e+17, 1.288743901648982e+17, 1.288743901688045e+17, 1.288743901728669e+17, 1.288743901767732e+17, 1.288743901808358e+17, 1.288743901848983e+17, 1.288743901888045e+17, 1.288743901928669e+17, 1.288743901967732e+17, 1.288743902008357e+17, 1.288743902048982e+17, 1.288743902088045e+17, 1.288743902128669e+17, 1.288743902167732e+17, 1.288743902208357e+17, 1.288743902248983e+17, 1.288743902288045e+17, 1.288743902328669e+17, 1.288743902367732e+17, 1.288743902408357e+17, 1.288743902448982e+17, 1.288743902488045e+17, 1.288743902528669e+17, 1.288743902567732e+17, 1.288743902608357e+17, 1.288743902648983e+17, 1.288743902688045e+17, 1.288743902728671e+17, 1.288743902767732e+17, 1.288743902808357e+17, 1.288743902848983e+17, 1.288743902888045e+17, 1.288743902928669e+17, 1.288743902967732e+17, 1.288743903008357e+17, 1.288743903048983e+17, 1.288743903088045e+17, 1.288743903128671e+17, 1.288743903167732e+17, 1.288743903208357e+17, 1.288743903248983e+17, 1.288743903288045e+17, 1.288743903328671e+17, 1.288743903367732e+17, 1.288743903408357e+17, 1.288743903448983e+17, 1.288743903488045e+17, 1.288743903528671e+17, 1.288743903567732e+17, 1.288743903608357e+17, 1.288743903648983e+17, 1.288743903688045e+17, 1.288743903728671e+17, 1.288743903767732e+17, 1.288743903808357e+17, 1.288743903848983e+17, 1.288743903888045e+17, 1.288743903928671e+17, 1.288743903967732e+17, 1.288743904008358e+17, 1.288743904048982e+17, 1.288743904088045e+17, 1.288743904128671e+17, 1.288743904167732e+17, 1.288743904208357e+17, 1.288743904248982e+17, 1.288743904288045e+17, 1.288743904328669e+17, 1.288743904367732e+17, 1.288743904408358e+17, 1.288743904448983e+17, 1.288743904488045e+17, 1.288743904528669e+17, 1.288743904567732e+17, 1.288743904608357e+17, 1.288743904648982e+17, 1.288743904688045e+17, 1.288743904728669e+17, 1.288743904767732e+17, 1.288743904808357e+17, 1.288743904848983e+17, 1.288743904888045e+17, 1.288743904928669e+17, 1.288743904967732e+17, 1.288743905008357e+17, 1.288743905048983e+17, 1.288743905088045e+17, 1.288743905128669e+17, 1.288743905167732e+17, 1.288743905208357e+17, 1.288743905248983e+17, 1.288743905288045e+17, 1.288743905328671e+17, 1.288743905367732e+17, 1.288743905408357e+17, 1.288743905448983e+17, 1.288743905488045e+17, 1.288743905528669e+17, 1.288743905567732e+17, 1.288743905608357e+17, 1.288743905648983e+17, 1.288743905688045e+17, 1.288743905728671e+17, 1.288743905767732e+17, 1.288743905808357e+17, 1.288743905848983e+17, 1.288743905888045e+17, 1.288743905928671e+17, 1.288743905967732e+17, 1.288743906008357e+17, 1.288743906048983e+17, 1.288743906088045e+17, 1.288743906128671e+17, 1.288743906167732e+17, 1.288743906208357e+17, 1.288743906248983e+17, 1.288743906288045e+17, 1.288743906328671e+17, 1.288743906367732e+17, 1.288743906408357e+17, 1.288743906448983e+17, 1.288743906488045e+17, 1.288743906528671e+17, 1.288743906567732e+17, 1.288743906608358e+17, 1.288743906648982e+17, 1.288743906688045e+17, 1.288743906728671e+17, 1.288743906767732e+17, 1.288743906808357e+17, 1.288743906848982e+17, 1.288743906888045e+17, 1.288743906928669e+17, 1.288743906967732e+17, 1.288743907008358e+17, 1.288743907048983e+17, 1.288743907088046e+17, 1.288743907128669e+17, 1.288743907167732e+17, 1.288743907208357e+17, 1.288743907248982e+17, 1.288743907288045e+17, 1.288743907328669e+17, 1.288743907367732e+17, 1.288743907408357e+17, 1.288743907448983e+17, 1.288743907488045e+17, 1.288743907528669e+17, 1.288743907567732e+17, 1.288743907608357e+17, 1.288743907648983e+17, 1.288743907688045e+17, 1.288743907728669e+17, 1.288743907767732e+17, 1.288743907808357e+17, 1.288743907848983e+17, 1.288743907888045e+17, 1.288743907928671e+17, 1.288743907967732e+17, 1.288743908008357e+17, 1.288743908048983e+17, 1.288743908088045e+17, 1.288743908128669e+17, 1.288743908167732e+17, 1.288743908208357e+17, 1.288743908248983e+17, 1.288743908288045e+17, 1.288743908328671e+17, 1.288743908367732e+17, 1.288743908408357e+17, 1.288743908448983e+17, 1.288743908488045e+17, 1.288743908528671e+17, 1.288743908567732e+17, 1.288743908608357e+17, 1.288743908648983e+17, 1.288743908688045e+17, 1.288743908728671e+17, 1.288743908767732e+17, 1.288743908808357e+17, 1.288743908848983e+17, 1.288743908888045e+17, 1.288743908928671e+17, 1.288743908967732e+17, 1.288743909008357e+17, 1.288743909048983e+17, 1.288743909088045e+17, 1.288743909128671e+17, 1.288743909167732e+17, 1.288743909208358e+17, 1.288743909248982e+17, 1.288743909288045e+17, 1.288743909328671e+17, 1.288743909367732e+17, 1.288743909408357e+17, 1.288743909448982e+17, 1.288743909488045e+17, 1.288743909528669e+17, 1.288743909567732e+17, 1.288743909608358e+17, 1.288743909648983e+17, 1.288743909688046e+17, 1.288743909728669e+17, 1.288743909767732e+17, 1.288743909808357e+17, 1.288743909848982e+17, 1.288743909888045e+17, 1.288743909928669e+17, 1.288743909967732e+17, 1.288743910008357e+17, 1.288743910048983e+17, 1.288743910088045e+17, 1.288743910128669e+17, 1.288743910167732e+17, 1.288743910208357e+17, 1.288743910248983e+17, 1.288743910288045e+17, 1.288743910328669e+17, 1.288743910367732e+17, 1.288743910408357e+17, 1.288743910448983e+17, 1.288743910488045e+17, 1.288743910528671e+17, 1.288743910567732e+17, 1.288743910608357e+17, 1.288743910648983e+17, 1.288743910688045e+17, 1.288743910728669e+17, 1.288743910767732e+17, 1.288743910808357e+17, 1.288743910848983e+17, 1.288743910888045e+17, 1.288743910928671e+17, 1.288743910967732e+17, 1.288743911008357e+17, 1.288743911048983e+17, 1.288743911088045e+17, 1.288743911128671e+17, 1.288743911167732e+17, 1.288743911208357e+17, 1.288743911248983e+17, 1.288743911288045e+17, 1.288743911328671e+17, 1.288743911367732e+17, 1.288743911408357e+17, 1.288743911448983e+17, 1.288743911488045e+17, 1.288743911528671e+17, 1.288743911567732e+17, 1.288743911608357e+17, 1.288743911648982e+17, 1.288743911688045e+17, 1.288743911728671e+17, 1.288743911767732e+17, 1.288743911808358e+17, 1.288743911848982e+17, 1.288743911888045e+17, 1.288743911928669e+17, 1.288743911967732e+17, 1.288743912008357e+17, 1.288743912048982e+17, 1.288743912088045e+17, 1.288743912128669e+17, 1.288743912167732e+17, 1.288743912208357e+17, 1.288743912248983e+17, 1.288743912288046e+17, 1.288743912328669e+17, 1.288743912367732e+17, 1.288743912408357e+17, 1.288743912448982e+17, 1.288743912488045e+17, 1.288743912528669e+17, 1.288743912567732e+17, 1.288743912608357e+17, 1.288743912648983e+17, 1.288743912688045e+17, 1.288743912728669e+17, 1.288743912767732e+17, 1.288743912808357e+17, 1.288743912848983e+17, 1.288743912888045e+17, 1.288743912928669e+17, 1.288743912967732e+17, 1.288743913008357e+17, 1.288743913048983e+17, 1.288743913088045e+17, 1.288743913128671e+17, 1.288743913167732e+17, 1.288743913208357e+17, 1.288743913248983e+17, 1.288743913288045e+17, 1.288743913328669e+17, 1.288743913367732e+17, 1.288743913408357e+17, 1.288743913448983e+17, 1.288743913488045e+17, 1.288743913528671e+17, 1.288743913567732e+17, 1.288743913608357e+17, 1.288743913648983e+17, 1.288743913688045e+17, 1.288743913728671e+17, 1.288743913767732e+17, 1.288743913808357e+17, 1.288743913848983e+17, 1.288743913888045e+17, 1.288743913928671e+17, 1.288743913967732e+17, 1.288743914008358e+17, 1.288743914048983e+17, 1.288743914088045e+17, 1.288743914128671e+17, 1.288743914167732e+17, 1.288743914208357e+17, 1.288743914248982e+17, 1.288743914288045e+17, 1.288743914328671e+17, 1.288743914367732e+17, 1.288743914408358e+17, 1.288743914448982e+17, 1.288743914488045e+17, 1.288743914528669e+17, 1.288743914567732e+17, 1.288743914608357e+17, 1.288743914648982e+17, 1.288743914688045e+17, 1.288743914728669e+17, 1.288743914767732e+17, 1.288743914808357e+17, 1.288743914848983e+17, 1.288743914888046e+17, 1.288743914928669e+17, 1.288743914967732e+17, 1.288743915008357e+17, 1.288743915048982e+17, 1.288743915088045e+17, 1.288743915128669e+17, 1.288743915167732e+17, 1.288743915208357e+17, 1.288743915248983e+17, 1.288743915288045e+17, 1.288743915328671e+17, 1.288743915367732e+17, 1.288743915408357e+17, 1.288743915448983e+17, 1.288743915488045e+17, 1.288743915528669e+17, 1.288743915567732e+17, 1.288743915608357e+17, 1.288743915648983e+17, 1.288743915688045e+17, 1.288743915728671e+17, 1.288743915767732e+17, 1.288743915808357e+17, 1.288743915848983e+17, 1.288743915888045e+17, 1.288743915928669e+17, 1.288743915967732e+17, 1.288743916008357e+17, 1.288743916048983e+17, 1.288743916088045e+17, 1.288743916128671e+17, 1.288743916167732e+17, 1.288743916208357e+17, 1.288743916248983e+17, 1.288743916288045e+17, 1.288743916328671e+17, 1.288743916367732e+17, 1.288743916408357e+17, 1.288743916448983e+17, 1.288743916488045e+17, 1.288743916528671e+17, 1.288743916567732e+17, 1.288743916608358e+17, 1.288743916648983e+17, 1.288743916688045e+17, 1.288743916728671e+17, 1.288743916767732e+17, 1.288743916808357e+17, 1.288743916848982e+17, 1.288743916888045e+17, 1.288743916928671e+17, 1.288743916967732e+17, 1.288743917008358e+17, 1.288743917048982e+17, 1.288743917088045e+17, 1.288743917128669e+17, 1.288743917167732e+17, 1.288743917208358e+17, 1.288743917248982e+17, 1.288743917288045e+17, 1.288743917328669e+17, 1.288743917367732e+17, 1.288743917408357e+17, 1.288743917448983e+17, 1.288743917488046e+17, 1.288743917528669e+17, 1.288743917567732e+17, 1.288743917608357e+17, 1.288743917648982e+17, 1.288743917688045e+17, 1.288743917728669e+17, 1.288743917767732e+17, 1.288743917808357e+17, 1.288743917848983e+17, 1.288743917888045e+17, 1.288743917928671e+17, 1.288743917967732e+17, 1.288743918008357e+17, 1.288743918048983e+17, 1.288743918088045e+17, 1.288743918128669e+17, 1.288743918167732e+17, 1.288743918208357e+17, 1.288743918248983e+17, 1.288743918288045e+17, 1.288743918328671e+17, 1.288743918367732e+17, 1.288743918408357e+17, 1.288743918448983e+17, 1.288743918488045e+17, 1.288743918528671e+17, 1.288743918567731e+17, 1.288743918608357e+17, 1.288743918648983e+17, 1.288743918688045e+17, 1.288743918728671e+17, 1.288743918767732e+17, 1.288743918808357e+17, 1.288743918848983e+17, 1.288743918888045e+17, 1.288743918928671e+17, 1.288743918967732e+17, 1.288743919008357e+17, 1.288743919048983e+17, 1.288743919088045e+17, 1.288743919128671e+17, 1.288743919167732e+17, 1.288743919208358e+17, 1.288743919248983e+17, 1.288743919288045e+17, 1.288743919328671e+17, 1.288743919367732e+17, 1.288743919408357e+17, 1.288743919448982e+17, 1.288743919488045e+17, 1.288743919528671e+17, 1.288743919567732e+17, 1.288743919608358e+17, 1.288743919648982e+17, 1.288743919688045e+17, 1.288743919728669e+17, 1.288743919767732e+17, 1.288743919808358e+17, 1.288743919848982e+17, 1.288743919888045e+17, 1.288743919928669e+17, 1.288743919967732e+17, 1.288743920008357e+17, 1.288743920048983e+17, 1.288743920088046e+17, 1.288743920128669e+17, 1.288743920167732e+17, 1.288743920208357e+17, 1.288743920248982e+17, 1.288743920288045e+17, 1.288743920328669e+17, 1.288743920367732e+17, 1.288743920408357e+17, 1.288743920448983e+17, 1.288743920488045e+17, 1.288743920528671e+17, 1.288743920567732e+17, 1.288743920608357e+17, 1.288743920648983e+17, 1.288743920688045e+17, 1.288743920728669e+17, 1.288743920767732e+17, 1.288743920808357e+17, 1.288743920848983e+17, 1.288743920888045e+17, 1.288743920928671e+17, 1.288743920967732e+17, 1.288743921008357e+17, 1.288743921048983e+17, 1.288743921088045e+17, 1.288743921128671e+17, 1.288743921167731e+17, 1.288743921208357e+17, 1.288743921248983e+17, 1.288743921288045e+17, 1.288743921328671e+17, 1.288743921367732e+17, 1.288743921408357e+17, 1.288743921448983e+17, 1.288743921488045e+17, 1.288743921528671e+17, 1.288743921567732e+17, 1.288743921608357e+17, 1.288743921648983e+17, 1.288743921688045e+17, 1.288743921728671e+17, 1.288743921767732e+17, 1.288743921808358e+17, 1.288743921848982e+17, 1.288743921888045e+17, 1.288743921928671e+17, 1.288743921967732e+17, 1.288743922008357e+17, 1.288743922048982e+17, 1.288743922088045e+17, 1.288743922128669e+17, 1.288743922167732e+17, 1.288743922208358e+17, 1.288743922248983e+17, 1.288743922288045e+17, 1.288743922328669e+17, 1.288743922367732e+17, 1.288743922408357e+17, 1.288743922448982e+17, 1.288743922488045e+17, 1.288743922528669e+17, 1.288743922567732e+17, 1.288743922608357e+17, 1.288743922648983e+17, 1.288743922688045e+17, 1.288743922728669e+17, 1.288743922767732e+17, 1.288743922808357e+17, 1.288743922848983e+17, 1.288743922888045e+17, 1.288743922928669e+17, 1.288743922967732e+17, 1.288743923008357e+17, 1.288743923048983e+17, 1.288743923088045e+17, 1.288743923128671e+17, 1.288743923167732e+17, 1.288743923208357e+17, 1.288743923248983e+17, 1.288743923288045e+17, 1.288743923328669e+17, 1.288743923367732e+17, 1.288743923408357e+17, 1.288743923448983e+17, 1.288743923488045e+17, 1.288743923528671e+17, 1.288743923567732e+17, 1.288743923608357e+17, 1.288743923648983e+17, 1.288743923688045e+17, 1.288743923728671e+17, 1.288743923767732e+17, 1.288743923808357e+17, 1.288743923848983e+17, 1.288743923888045e+17, 1.288743923928671e+17, 1.288743923967732e+17, 1.288743924008357e+17, 1.288743924048983e+17, 1.288743924088045e+17, 1.288743924128671e+17, 1.288743924167732e+17, 1.288743924208357e+17, 1.288743924248983e+17, 1.288743924288045e+17, 1.288743924328671e+17, 1.288743924367732e+17, 1.288743924408358e+17, 1.288743924448982e+17, 1.288743924488045e+17, 1.288743924528671e+17, 1.288743924567732e+17, 1.288743924608357e+17, 1.288743924648982e+17, 1.288743924688045e+17, 1.288743924728669e+17, 1.288743924767732e+17, 1.288743924808358e+17, 1.288743924848983e+17, 1.288743924888045e+17, 1.288743924928669e+17, 1.288743924967732e+17, 1.288743925008357e+17, 1.288743925048982e+17, 1.288743925088045e+17, 1.288743925128669e+17, 1.288743925167732e+17, 1.288743925208357e+17, 1.288743925248983e+17, 1.288743925288045e+17, 1.288743925328669e+17, 1.288743925367732e+17, 1.288743925408357e+17, 1.288743925448983e+17, 1.288743925488045e+17, 1.288743925528669e+17, 1.288743925567732e+17, 1.288743925608357e+17, 1.288743925648983e+17, 1.288743925688045e+17, 1.288743925728671e+17, 1.288743925767732e+17, 1.288743925808357e+17, 1.288743925848983e+17, 1.288743925888045e+17, 1.288743925928669e+17, 1.288743925967732e+17, 1.288743926008357e+17, 1.288743926048983e+17, 1.288743926088045e+17, 1.288743926128671e+17, 1.288743926167732e+17, 1.288743926208357e+17, 1.288743926248983e+17, 1.288743926288045e+17, 1.288743926328671e+17, 1.288743926367732e+17, 1.288743926408357e+17, 1.288743926448983e+17, 1.288743926488045e+17, 1.288743926528671e+17, 1.288743926567732e+17, 1.288743926608357e+17, 1.288743926648983e+17, 1.288743926688045e+17, 1.288743926728671e+17, 1.288743926767732e+17, 1.288743926808357e+17, 1.288743926848983e+17, 1.288743926888045e+17, 1.288743926928671e+17, 1.288743926967732e+17, 1.288743927008358e+17, 1.288743927048982e+17, 1.288743927088045e+17, 1.288743927128671e+17, 1.288743927167732e+17, 1.288743927208357e+17, 1.288743927248982e+17, 1.288743927288045e+17, 1.288743927328669e+17, 1.288743927367732e+17, 1.288743927408358e+17, 1.288743927448983e+17, 1.288743927488046e+17, 1.288743927528669e+17, 1.288743927567732e+17, 1.288743927608357e+17, 1.288743927648982e+17, 1.288743927688045e+17, 1.288743927728669e+17, 1.288743927767732e+17, 1.288743927808357e+17, 1.288743927848983e+17, 1.288743927888045e+17, 1.288743927928669e+17, 1.288743927967732e+17, 1.288743928008357e+17, 1.288743928048983e+17, 1.288743928088045e+17, 1.288743928128669e+17, 1.288743928167732e+17, 1.288743928208357e+17, 1.288743928248983e+17, 1.288743928288045e+17, 1.288743928328671e+17, 1.288743928367732e+17, 1.288743928408357e+17, 1.288743928448983e+17, 1.288743928488045e+17, 1.288743928528669e+17, 1.288743928567732e+17, 1.288743928608357e+17, 1.288743928648983e+17, 1.288743928688045e+17, 1.288743928728671e+17, 1.288743928767732e+17, 1.288743928808357e+17, 1.288743928848983e+17, 1.288743928888045e+17, 1.288743928928671e+17, 1.288743928967732e+17, 1.288743929008357e+17, 1.288743929048983e+17, 1.288743929088045e+17, 1.288743929128671e+17, 1.288743929167732e+17, 1.288743929208357e+17, 1.288743929248983e+17, 1.288743929288045e+17, 1.288743929328671e+17, 1.288743929367732e+17, 1.288743929408357e+17, 1.288743929448983e+17, 1.288743929488045e+17, 1.288743929528671e+17, 1.288743929567732e+17, 1.288743929608358e+17, 1.288743929648982e+17, 1.288743929688045e+17, 1.288743929728671e+17, 1.288743929767732e+17, 1.288743929808357e+17, 1.288743929848982e+17, 1.288743929888045e+17, 1.288743929928669e+17, 1.288743929967732e+17, 1.288743930008358e+17, 1.288743930048983e+17, 1.288743930088046e+17, 1.288743930128669e+17, 1.288743930167732e+17, 1.288743930208357e+17, 1.288743930248982e+17, 1.288743930288045e+17, 1.288743930328669e+17, 1.288743930367732e+17, 1.288743930408357e+17, 1.288743930448983e+17, 1.288743930488045e+17, 1.288743930528669e+17, 1.288743930567732e+17, 1.288743930608357e+17, 1.288743930648983e+17, 1.288743930688045e+17, 1.288743930728669e+17, 1.288743930767732e+17, 1.288743930808357e+17, 1.288743930848983e+17, 1.288743930888045e+17, 1.288743930928671e+17, 1.288743930967732e+17, 1.288743931008357e+17, 1.288743931048983e+17, 1.288743931088045e+17, 1.288743931128669e+17, 1.288743931167732e+17, 1.288743931208357e+17, 1.288743931248983e+17, 1.288743931288045e+17, 1.288743931328671e+17, 1.288743931367732e+17, 1.288743931408357e+17, 1.288743931448983e+17, 1.288743931488045e+17, 1.288743931528671e+17, 1.288743931567732e+17, 1.288743931608357e+17, 1.288743931648983e+17, 1.288743931688045e+17, 1.288743931728671e+17, 1.288743931767732e+17, 1.288743931808357e+17, 1.288743931848983e+17, 1.288743931888045e+17, 1.288743931928671e+17, 1.288743931967732e+17, 1.288743932008357e+17, 1.288743932048982e+17, 1.288743932088045e+17, 1.288743932128671e+17, 1.288743932167732e+17, 1.288743932208358e+17, 1.288743932248982e+17, 1.288743932288045e+17, 1.288743932328669e+17, 1.288743932367732e+17, 1.288743932408357e+17, 1.288743932448982e+17, 1.288743932488045e+17, 1.288743932528669e+17, 1.288743932567732e+17, 1.288743932608357e+17, 1.288743932648983e+17, 1.288743932688046e+17, 1.288743932728669e+17, 1.288743932767732e+17, 1.288743932808357e+17, 1.288743932848982e+17, 1.288743932888045e+17, 1.288743932928669e+17, 1.288743932967732e+17, 1.288743933008357e+17, 1.288743933048983e+17, 1.288743933088045e+17, 1.288743933128669e+17, 1.288743933167732e+17, 1.288743933208357e+17, 1.288743933248983e+17, 1.288743933288045e+17, 1.288743933328669e+17, 1.288743933367732e+17, 1.288743933408357e+17, 1.288743933448983e+17, 1.288743933488045e+17, 1.288743933528671e+17, 1.288743933567732e+17, 1.288743933608357e+17, 1.288743933648983e+17, 1.288743933688045e+17, 1.288743933728669e+17, 1.288743933767732e+17, 1.288743933808357e+17, 1.288743933848983e+17, 1.288743933888045e+17, 1.288743933928671e+17, 1.288743933967732e+17, 1.288743934008357e+17, 1.288743934048983e+17, 1.288743934088045e+17, 1.288743934128671e+17, 1.288743934167732e+17, 1.288743934208357e+17, 1.288743934248983e+17, 1.288743934288045e+17, 1.288743934328671e+17, 1.288743934367732e+17, 1.288743934408358e+17, 1.288743934448983e+17, 1.288743934488045e+17, 1.288743934528671e+17, 1.288743934567732e+17, 1.288743934608357e+17, 1.288743934648982e+17, 1.288743934688045e+17, 1.288743934728671e+17, 1.288743934767732e+17, 1.288743934808358e+17, 1.288743934848982e+17, 1.288743934888045e+17, 1.288743934928669e+17, 1.288743934967732e+17, 1.288743935008358e+17, 1.288743935048982e+17, 1.288743935088045e+17, 1.288743935128669e+17, 1.288743935167732e+17, 1.288743935208357e+17, 1.288743935248983e+17, 1.288743935288046e+17, 1.288743935328669e+17, 1.288743935367732e+17, 1.288743935408357e+17, 1.288743935448982e+17, 1.288743935488045e+17, 1.288743935528669e+17, 1.288743935567732e+17, 1.288743935608357e+17, 1.288743935648983e+17, 1.288743935688045e+17, 1.288743935728671e+17, 1.288743935767732e+17, 1.288743935808357e+17, 1.288743935848983e+17, 1.288743935888045e+17, 1.288743935928669e+17, 1.288743935967732e+17, 1.288743936008357e+17, 1.288743936048983e+17, 1.288743936088045e+17, 1.288743936128671e+17, 1.288743936167732e+17, 1.288743936208357e+17, 1.288743936248983e+17, 1.288743936288045e+17, 1.288743936328671e+17, 1.288743936367731e+17, 1.288743936408357e+17, 1.288743936448983e+17, 1.288743936488045e+17, 1.288743936528671e+17, 1.288743936567732e+17, 1.288743936608357e+17, 1.288743936648983e+17, 1.288743936688045e+17, 1.288743936728671e+17, 1.288743936767732e+17, 1.288743936808357e+17, 1.288743936848983e+17, 1.288743936888045e+17, 1.288743936928671e+17, 1.288743936967732e+17, 1.288743937008358e+17, 1.288743937048983e+17, 1.288743937088045e+17, 1.288743937128671e+17, 1.288743937167732e+17, 1.288743937208357e+17, 1.288743937248982e+17, 1.288743937288045e+17, 1.288743937328671e+17, 1.288743937367732e+17, 1.288743937408358e+17, 1.288743937448982e+17, 1.288743937488045e+17, 1.288743937528669e+17, 1.288743937567732e+17, 1.288743937608358e+17, 1.288743937648982e+17, 1.288743937688045e+17, 1.288743937728669e+17, 1.288743937767732e+17, 1.288743937808357e+17, 1.288743937848983e+17, 1.288743937888046e+17, 1.288743937928669e+17, 1.288743937967732e+17, 1.288743938008357e+17, 1.288743938048982e+17, 1.288743938088045e+17, 1.288743938128669e+17, 1.288743938167732e+17, 1.288743938208357e+17, 1.288743938248983e+17, 1.288743938288045e+17, 1.288743938328671e+17, 1.288743938367732e+17, 1.288743938408357e+17, 1.288743938448983e+17, 1.288743938488045e+17, 1.288743938528669e+17, 1.288743938567732e+17, 1.288743938608357e+17, 1.288743938648983e+17, 1.288743938688045e+17, 1.288743938728671e+17, 1.288743938767732e+17, 1.288743938808357e+17, 1.288743938848983e+17, 1.288743938888045e+17, 1.288743938928671e+17, 1.288743938967731e+17, 1.288743939008357e+17, 1.288743939048983e+17, 1.288743939088045e+17, 1.288743939128671e+17, 1.288743939167732e+17, 1.288743939208357e+17, 1.288743939248983e+17, 1.288743939288045e+17, 1.288743939328671e+17, 1.288743939367732e+17, 1.288743939408357e+17, 1.288743939448983e+17, 1.288743939488045e+17, 1.288743939528671e+17, 1.288743939567732e+17, 1.288743939608358e+17, 1.288743939648982e+17, 1.288743939688045e+17, 1.288743939728671e+17, 1.288743939767732e+17, 1.288743939808357e+17, 1.288743939848982e+17, 1.288743939888045e+17, 1.288743939928669e+17, 1.288743939967732e+17, 1.288743940008358e+17, 1.288743940048983e+17, 1.288743940088045e+17, 1.288743940128669e+17, 1.288743940167732e+17, 1.288743940208357e+17, 1.288743940248982e+17, 1.288743940288045e+17, 1.288743940328669e+17, 1.288743940367732e+17, 1.288743940408357e+17, 1.288743940448983e+17, 1.288743940488045e+17, 1.288743940528669e+17, 1.288743940567732e+17, 1.288743940608357e+17, 1.288743940648982e+17, 1.288743940688045e+17, 1.288743940728669e+17, 1.288743940767732e+17, 1.288743940808357e+17, 1.288743940848983e+17, 1.288743940888045e+17, 1.288743940928671e+17, 1.288743940967732e+17, 1.288743941008357e+17, 1.288743941048983e+17, 1.288743941088045e+17, 1.288743941128669e+17, 1.288743941167732e+17, 1.288743941208357e+17, 1.288743941248983e+17, 1.288743941288045e+17, 1.288743941328671e+17, 1.288743941367732e+17, 1.288743941408357e+17, 1.288743941448983e+17, 1.288743941488045e+17, 1.288743941528671e+17, 1.288743941567732e+17, 1.288743941608357e+17, 1.288743941648983e+17, 1.288743941688045e+17, 1.288743941728671e+17, 1.288743941767732e+17, 1.288743941808357e+17, 1.288743941848983e+17, 1.288743941888045e+17, 1.288743941928671e+17, 1.288743941967732e+17, 1.288743942008357e+17, 1.288743942048983e+17, 1.288743942088045e+17, 1.288743942128671e+17, 1.288743942167732e+17, 1.288743942208358e+17, 1.288743942248982e+17, 1.288743942288045e+17, 1.288743942328671e+17, 1.288743942367732e+17, 1.288743942408357e+17, 1.288743942448982e+17, 1.288743942488045e+17, 1.288743942528669e+17, 1.288743942567732e+17, 1.288743942608358e+17, 1.288743942648983e+17, 1.288743942688045e+17, 1.288743942728669e+17, 1.288743942767732e+17, 1.288743942808357e+17, 1.288743942848982e+17, 1.288743942888045e+17, 1.288743942928669e+17, 1.288743942967732e+17, 1.288743943008357e+17, 1.288743943048983e+17, 1.288743943088045e+17, 1.288743943128669e+17, 1.288743943167732e+17, 1.288743943208357e+17, 1.288743943248983e+17, 1.288743943288045e+17, 1.288743943328669e+17, 1.288743943367732e+17, 1.288743943408357e+17, 1.288743943448983e+17, 1.288743943488045e+17, 1.288743943528671e+17, 1.288743943567732e+17, 1.288743943608357e+17, 1.288743943648983e+17, 1.288743943688045e+17, 1.288743943728669e+17, 1.288743943767732e+17, 1.288743943808357e+17, 1.288743943848983e+17, 1.288743943888045e+17, 1.288743943928671e+17, 1.288743943967732e+17, 1.288743944008357e+17, 1.288743944048983e+17, 1.288743944088045e+17, 1.288743944128671e+17, 1.288743944167732e+17, 1.288743944208357e+17, 1.288743944248983e+17, 1.288743944288045e+17, 1.288743944328671e+17, 1.288743944367732e+17, 1.288743944408357e+17, 1.288743944448983e+17, 1.288743944488045e+17, 1.288743944528671e+17, 1.288743944567732e+17, 1.288743944608357e+17, 1.288743944648983e+17, 1.288743944688045e+17, 1.288743944728671e+17, 1.288743944767732e+17, 1.288743944808358e+17, 1.288743944848982e+17, 1.288743944888045e+17, 1.288743944928671e+17, 1.288743944967732e+17, 1.288743945008357e+17, 1.288743945048982e+17, 1.288743945088045e+17, 1.288743945128669e+17, 1.288743945167732e+17, 1.288743945208358e+17, 1.288743945248983e+17, 1.288743945288046e+17, 1.288743945328669e+17, 1.288743945367732e+17, 1.288743945408357e+17, 1.288743945448982e+17, 1.288743945488045e+17, 1.288743945528669e+17, 1.288743945567732e+17, 1.288743945608357e+17, 1.288743945648983e+17, 1.288743945688045e+17, 1.288743945728669e+17, 1.288743945767732e+17, 1.288743945808357e+17, 1.288743945848983e+17, 1.288743945888045e+17, 1.288743945928669e+17, 1.288743945967732e+17, 1.288743946008357e+17, 1.288743946048983e+17, 1.288743946088045e+17, 1.288743946128671e+17, 1.288743946167732e+17, 1.288743946208357e+17, 1.288743946248983e+17, 1.288743946288045e+17, 1.288743946328669e+17, 1.288743946367732e+17, 1.288743946408357e+17, 1.288743946448983e+17, 1.288743946488045e+17, 1.288743946528671e+17, 1.288743946567732e+17, 1.288743946608357e+17, 1.288743946648983e+17, 1.288743946688045e+17, 1.288743946728671e+17, 1.288743946767732e+17, 1.288743946808357e+17, 1.288743946848983e+17, 1.288743946888045e+17, 1.288743946928671e+17, 1.288743946967732e+17, 1.288743947008357e+17, 1.288743947048983e+17, 1.288743947088045e+17, 1.288743947128671e+17, 1.288743947167732e+17, 1.288743947208357e+17, 1.288743947248983e+17, 1.288743947288045e+17, 1.288743947328671e+17, 1.288743947367732e+17, 1.288743947408358e+17, 1.288743947448982e+17, 1.288743947488045e+17, 1.288743947528671e+17, 1.288743947567732e+17, 1.288743947608357e+17, 1.288743947648982e+17, 1.288743947688045e+17, 1.288743947728669e+17, 1.288743947767732e+17, 1.288743947808358e+17, 1.288743947848983e+17, 1.288743947888046e+17, 1.288743947928669e+17, 1.288743947967732e+17, 1.288743948008357e+17, 1.288743948048982e+17, 1.288743948088045e+17, 1.288743948128669e+17, 1.288743948167732e+17, 1.288743948208357e+17, 1.288743948248983e+17, 1.288743948288045e+17, 1.288743948328669e+17, 1.288743948367732e+17, 1.288743948408357e+17, 1.288743948448983e+17, 1.288743948488045e+17, 1.288743948528669e+17, 1.288743948567732e+17, 1.288743948608357e+17, 1.288743948648983e+17, 1.288743948688045e+17, 1.288743948728671e+17, 1.288743948767732e+17, 1.288743948808357e+17, 1.288743948848983e+17, 1.288743948888045e+17, 1.288743948928669e+17, 1.288743948967732e+17, 1.288743949008357e+17, 1.288743949048983e+17, 1.288743949088045e+17, 1.288743949128671e+17, 1.288743949167732e+17, 1.288743949208357e+17, 1.288743949248983e+17, 1.288743949288045e+17, 1.288743949328671e+17, 1.288743949367732e+17, 1.288743949408357e+17, 1.288743949448983e+17, 1.288743949488045e+17, 1.288743949528671e+17, 1.288743949567732e+17, 1.288743949608357e+17, 1.288743949648983e+17, 1.288743949688045e+17, 1.288743949728671e+17, 1.288743949767732e+17, 1.288743949808357e+17, 1.288743949848982e+17, 1.288743949888045e+17, 1.288743949928671e+17, 1.288743949967732e+17, 1.288743950008358e+17, 1.288743950048982e+17, 1.288743950088045e+17, 1.288743950128669e+17, 1.288743950167732e+17, 1.288743950208357e+17, 1.288743950248982e+17, 1.288743950288045e+17, 1.288743950328669e+17, 1.288743950367732e+17, 1.288743950408357e+17, 1.288743950448983e+17, 1.288743950488046e+17, 1.288743950528669e+17, 1.288743950567732e+17, 1.288743950608357e+17, 1.288743950648982e+17, 1.288743950688045e+17, 1.288743950728669e+17, 1.288743950767732e+17, 1.288743950808357e+17, 1.288743950848983e+17, 1.288743950888045e+17, 1.288743950928669e+17, 1.288743950967732e+17, 1.288743951008357e+17, 1.288743951048983e+17, 1.288743951088045e+17, 1.288743951128669e+17, 1.288743951167732e+17, 1.288743951208357e+17, 1.288743951248983e+17, 1.288743951288045e+17, 1.288743951328671e+17, 1.288743951367732e+17, 1.288743951408357e+17, 1.288743951448983e+17, 1.288743951488045e+17, 1.288743951528669e+17, 1.288743951567732e+17, 1.288743951608357e+17, 1.288743951648983e+17, 1.288743951688045e+17, 1.288743951728671e+17, 1.288743951767732e+17, 1.288743951808357e+17, 1.288743951848983e+17, 1.288743951888045e+17, 1.288743951928671e+17, 1.288743951967732e+17, 1.288743952008357e+17, 1.288743952048983e+17, 1.288743952088045e+17, 1.288743952128671e+17, 1.288743952167732e+17, 1.288743952208358e+17, 1.288743952248983e+17, 1.288743952288045e+17, 1.288743952328671e+17, 1.288743952367732e+17, 1.288743952408357e+17, 1.288743952448982e+17, 1.288743952488045e+17, 1.288743952528671e+17, 1.288743952567732e+17, 1.288743952608358e+17, 1.288743952648982e+17, 1.288743952688045e+17, 1.288743952728669e+17, 1.288743952767732e+17, 1.288743952808357e+17, 1.288743952848982e+17, 1.288743952888045e+17, 1.288743952928669e+17, 1.288743952967732e+17, 1.288743953008357e+17, 1.288743953048983e+17, 1.288743953088046e+17, 1.288743953128669e+17, 1.288743953167732e+17, 1.288743953208357e+17, 1.288743953248982e+17, 1.288743953288045e+17, 1.288743953328669e+17, 1.288743953367732e+17, 1.288743953408357e+17, 1.288743953448983e+17, 1.288743953488045e+17, 1.288743953528671e+17, 1.288743953567732e+17, 1.288743953608357e+17, 1.288743953648983e+17, 1.288743953688045e+17, 1.288743953728669e+17, 1.288743953767732e+17, 1.288743953808357e+17, 1.288743953848983e+17, 1.288743953888045e+17, 1.288743953928671e+17, 1.288743953967732e+17, 1.288743954008357e+17, 1.288743954048983e+17, 1.288743954088045e+17, 1.288743954128669e+17, 1.288743954167732e+17, 1.288743954208357e+17, 1.288743954248983e+17, 1.288743954288045e+17, 1.288743954328671e+17, 1.288743954367732e+17, 1.288743954408357e+17, 1.288743954448983e+17, 1.288743954488045e+17, 1.288743954528671e+17, 1.288743954567732e+17, 1.288743954608357e+17, 1.288743954648983e+17, 1.288743954688045e+17, 1.288743954728671e+17, 1.288743954767732e+17, 1.288743954808358e+17, 1.288743954848983e+17, 1.288743954888045e+17, 1.288743954928671e+17, 1.288743954967732e+17, 1.288743955008357e+17, 1.288743955048982e+17, 1.288743955088045e+17, 1.288743955128671e+17, 1.288743955167732e+17, 1.288743955208358e+17, 1.288743955248982e+17, 1.288743955288045e+17, 1.288743955328669e+17, 1.288743955367732e+17, 1.288743955408358e+17, 1.288743955448982e+17, 1.288743955488045e+17, 1.288743955528669e+17, 1.288743955567732e+17, 1.288743955608357e+17, 1.288743955648983e+17, 1.288743955688046e+17, 1.288743955728669e+17, 1.288743955767732e+17, 1.288743955808357e+17, 1.288743955848982e+17, 1.288743955888045e+17, 1.288743955928669e+17, 1.288743955967732e+17, 1.288743956008357e+17, 1.288743956048983e+17, 1.288743956088045e+17, 1.288743956128671e+17, 1.288743956167732e+17, 1.288743956208357e+17, 1.288743956248983e+17, 1.288743956288045e+17, 1.288743956328669e+17, 1.288743956367732e+17, 1.288743956408357e+17, 1.288743956448983e+17, 1.288743956488045e+17, 1.288743956528671e+17, 1.288743956567732e+17, 1.288743956608357e+17, 1.288743956648983e+17, 1.288743956688045e+17, 1.288743956728671e+17, 1.288743956767731e+17, 1.288743956808357e+17, 1.288743956848983e+17, 1.288743956888045e+17, 1.288743956928671e+17, 1.288743956967732e+17, 1.288743957008357e+17, 1.288743957048983e+17, 1.288743957088045e+17, 1.288743957128671e+17, 1.288743957167732e+17, 1.288743957208357e+17, 1.288743957248983e+17, 1.288743957288045e+17, 1.288743957328671e+17, 1.288743957367732e+17, 1.288743957408358e+17, 1.288743957448983e+17, 1.288743957488045e+17, 1.288743957528671e+17, 1.288743957567732e+17, 1.288743957608357e+17, 1.288743957648982e+17, 1.288743957688045e+17, 1.288743957728671e+17, 1.288743957767732e+17, 1.288743957808358e+17, 1.288743957848982e+17, 1.288743957888045e+17, 1.288743957928669e+17, 1.288743957967732e+17, 1.288743958008358e+17, 1.288743958048982e+17, 1.288743958088045e+17, 1.288743958128669e+17, 1.288743958167732e+17, 1.288743958208357e+17, 1.288743958248983e+17, 1.288743958288046e+17, 1.288743958328669e+17, 1.288743958367732e+17, 1.288743958408357e+17, 1.288743958448982e+17, 1.288743958488045e+17, 1.288743958528669e+17, 1.288743958567732e+17, 1.288743958608357e+17, 1.288743958648983e+17, 1.288743958688045e+17, 1.288743958728671e+17, 1.288743958767732e+17, 1.288743958808357e+17, 1.288743958848983e+17, 1.288743958888045e+17, 1.288743958928669e+17, 1.288743958967732e+17, 1.288743959008357e+17, 1.288743959048983e+17, 1.288743959088045e+17, 1.288743959128671e+17, 1.288743959167732e+17, 1.288743959208357e+17, 1.288743959248983e+17, 1.288743959288045e+17, 1.288743959328671e+17, 1.288743959367731e+17, 1.288743959408357e+17, 1.288743959448983e+17, 1.288743959488045e+17, 1.288743959528671e+17, 1.288743959567732e+17, 1.288743959608357e+17, 1.288743959648983e+17, 1.288743959688045e+17, 1.288743959728671e+17, 1.288743959767732e+17, 1.288743959808357e+17, 1.288743959848983e+17, 1.288743959888045e+17, 1.288743959928671e+17, 1.288743959967732e+17, 1.288743960008358e+17, 1.288743960048982e+17, 1.288743960088045e+17, 1.288743960128671e+17, 1.288743960167732e+17, 1.288743960208357e+17, 1.288743960248982e+17, 1.288743960288045e+17, 1.288743960328669e+17, 1.288743960367732e+17, 1.288743960408358e+17, 1.288743960448983e+17, 1.288743960488045e+17, 1.288743960528669e+17, 1.288743960567732e+17, 1.288743960608357e+17, 1.288743960648982e+17, 1.288743960688045e+17, 1.288743960728669e+17, 1.288743960767732e+17, 1.288743960808357e+17, 1.288743960848983e+17, 1.288743960888045e+17, 1.288743960928669e+17, 1.288743960967732e+17, 1.288743961008357e+17, 1.288743961048982e+17, 1.288743961088045e+17, 1.288743961128669e+17, 1.288743961167732e+17, 1.288743961208357e+17, 1.288743961248983e+17, 1.288743961288045e+17, 1.288743961328671e+17, 1.288743961367732e+17, 1.288743961408357e+17, 1.288743961448983e+17, 1.288743961488045e+17, 1.288743961528669e+17, 1.288743961567732e+17, 1.288743961608357e+17, 1.288743961648983e+17, 1.288743961688045e+17, 1.288743961728671e+17, 1.288743961767732e+17, 1.288743961808357e+17, 1.288743961848983e+17, 1.288743961888045e+17, 1.288743961928671e+17, 1.288743961967732e+17, 1.288743962008357e+17, 1.288743962048983e+17, 1.288743962088045e+17, 1.288743962128671e+17, 1.288743962167732e+17, 1.288743962208357e+17, 1.288743962248983e+17, 1.288743962288045e+17, 1.288743962328671e+17, 1.288743962367732e+17, 1.288743962408357e+17, 1.288743962448983e+17, 1.288743962488045e+17, 1.288743962528671e+17, 1.288743962567732e+17, 1.288743962608358e+17, 1.288743962648982e+17, 1.288743962688045e+17, 1.288743962728671e+17, 1.288743962767732e+17, 1.288743962808357e+17, 1.288743962848982e+17, 1.288743962888045e+17, 1.288743962928669e+17, 1.288743962967732e+17, 1.288743963008358e+17, 1.288743963048983e+17, 1.288743963088045e+17, 1.288743963128669e+17, 1.288743963167732e+17, 1.288743963208357e+17, 1.288743963248982e+17, 1.288743963288045e+17, 1.288743963328669e+17, 1.288743963367732e+17, 1.288743963408357e+17, 1.288743963448983e+17, 1.288743963488045e+17, 1.288743963528669e+17, 1.288743963567732e+17, 1.288743963608357e+17, 1.288743963648983e+17, 1.288743963688045e+17, 1.288743963728669e+17, 1.288743963767732e+17, 1.288743963808357e+17, 1.288743963848983e+17, 1.288743963888045e+17, 1.288743963928671e+17, 1.288743963967732e+17, 1.288743964008357e+17, 1.288743964048983e+17, 1.288743964088045e+17, 1.288743964128669e+17, 1.288743964167732e+17, 1.288743964208357e+17, 1.288743964248983e+17, 1.288743964288045e+17, 1.288743964328671e+17, 1.288743964367732e+17, 1.288743964408357e+17, 1.288743964448983e+17, 1.288743964488045e+17, 1.288743964528671e+17, 1.288743964567732e+17, 1.288743964608357e+17, 1.288743964648983e+17, 1.288743964688045e+17, 1.288743964728671e+17, 1.288743964767732e+17, 1.288743964808357e+17, 1.288743964848983e+17, 1.288743964888045e+17, 1.288743964928671e+17, 1.288743964967732e+17, 1.288743965008357e+17, 1.288743965048983e+17, 1.288743965088045e+17, 1.288743965128671e+17, 1.288743965167732e+17, 1.288743965208358e+17, 1.288743965248982e+17, 1.288743965288045e+17, 1.288743965328671e+17, 1.288743965367732e+17, 1.288743965408357e+17, 1.288743965448982e+17, 1.288743965488045e+17, 1.288743965528669e+17, 1.288743965567732e+17, 1.288743965608358e+17, 1.288743965648983e+17, 1.288743965688046e+17, 1.288743965728669e+17, 1.288743965767732e+17, 1.288743965808357e+17, 1.288743965848982e+17, 1.288743965888045e+17, 1.288743965928669e+17, 1.288743965967732e+17, 1.288743966008357e+17, 1.288743966048983e+17, 1.288743966088045e+17, 1.288743966128669e+17, 1.288743966167732e+17, 1.288743966208357e+17, 1.288743966248983e+17, 1.288743966288045e+17, 1.288743966328669e+17, 1.288743966367732e+17, 1.288743966408357e+17, 1.288743966448983e+17, 1.288743966488045e+17, 1.288743966528671e+17, 1.288743966567732e+17, 1.288743966608357e+17, 1.288743966648983e+17, 1.288743966688045e+17, 1.288743966728669e+17, 1.288743966767732e+17, 1.288743966808357e+17, 1.288743966848983e+17, 1.288743966888045e+17, 1.288743966928671e+17, 1.288743966967732e+17, 1.288743967008357e+17, 1.288743967048983e+17, 1.288743967088045e+17, 1.288743967128671e+17, 1.288743967167732e+17, 1.288743967208357e+17, 1.288743967248983e+17, 1.288743967288045e+17, 1.288743967328671e+17, 1.288743967367732e+17, 1.288743967408357e+17, 1.288743967448983e+17, 1.288743967488045e+17, 1.288743967528671e+17, 1.288743967567732e+17, 1.288743967608357e+17, 1.288743967648983e+17, 1.288743967688045e+17, 1.288743967728671e+17, 1.288743967767732e+17, 1.288743967808358e+17, 1.288743967848982e+17, 1.288743967888045e+17, 1.288743967928671e+17, 1.288743967967732e+17, 1.288743968008357e+17, 1.288743968048982e+17, 1.288743968088045e+17, 1.288743968128669e+17, 1.288743968167732e+17, 1.288743968208358e+17, 1.288743968248983e+17, 1.288743968288046e+17, 1.288743968328669e+17, 1.288743968367732e+17, 1.288743968408357e+17, 1.288743968448982e+17, 1.288743968488045e+17, 1.288743968528669e+17, 1.288743968567732e+17, 1.288743968608357e+17, 1.288743968648983e+17, 1.288743968688045e+17, 1.288743968728669e+17, 1.288743968767732e+17, 1.288743968808357e+17, 1.288743968848983e+17, 1.288743968888045e+17, 1.288743968928669e+17, 1.288743968967732e+17, 1.288743969008357e+17, 1.288743969048983e+17, 1.288743969088045e+17, 1.288743969128671e+17, 1.288743969167732e+17, 1.288743969208357e+17, 1.288743969248983e+17, 1.288743969288045e+17, 1.288743969328669e+17, 1.288743969367732e+17, 1.288743969408357e+17, 1.288743969448983e+17, 1.288743969488045e+17, 1.288743969528671e+17, 1.288743969567732e+17, 1.288743969608357e+17, 1.288743969648983e+17, 1.288743969688045e+17, 1.288743969728671e+17, 1.288743969767732e+17, 1.288743969808357e+17, 1.288743969848983e+17, 1.288743969888045e+17, 1.288743969928671e+17, 1.288743969967732e+17, 1.288743970008357e+17, 1.288743970048983e+17, 1.288743970088045e+17, 1.288743970128671e+17, 1.288743970167732e+17, 1.288743970208357e+17, 1.288743970248982e+17, 1.288743970288045e+17, 1.288743970328671e+17, 1.288743970367732e+17, 1.288743970408358e+17, 1.288743970448982e+17, 1.288743970488045e+17, 1.288743970528669e+17, 1.288743970567732e+17, 1.288743970608357e+17, 1.288743970648982e+17, 1.288743970688045e+17, 1.288743970728669e+17, 1.288743970767732e+17, 1.288743970808357e+17, 1.288743970848983e+17, 1.288743970888046e+17, 1.288743970928669e+17, 1.288743970967732e+17, 1.288743971008357e+17, 1.288743971048982e+17, 1.288743971088045e+17, 1.288743971128669e+17, 1.288743971167732e+17, 1.288743971208357e+17, 1.288743971248983e+17, 1.288743971288045e+17, 1.288743971328669e+17, 1.288743971367732e+17, 1.288743971408357e+17, 1.288743971448983e+17, 1.288743971488045e+17, 1.288743971528669e+17, 1.288743971567732e+17, 1.288743971608357e+17, 1.288743971648983e+17, 1.288743971688045e+17, 1.288743971728671e+17, 1.288743971767732e+17, 1.288743971808357e+17, 1.288743971848983e+17, 1.288743971888045e+17, 1.288743971928669e+17, 1.288743971967732e+17, 1.288743972008357e+17, 1.288743972048983e+17, 1.288743972088045e+17, 1.288743972128671e+17, 1.288743972167732e+17, 1.288743972208357e+17, 1.288743972248983e+17, 1.288743972288045e+17, 1.288743972328671e+17, 1.288743972367732e+17, 1.288743972408357e+17, 1.288743972448983e+17, 1.288743972488045e+17, 1.288743972528671e+17, 1.288743972567732e+17, 1.288743972608358e+17, 1.288743972648983e+17, 1.288743972688045e+17, 1.288743972728671e+17, 1.288743972767732e+17, 1.288743972808357e+17, 1.288743972848982e+17, 1.288743972888045e+17, 1.288743972928671e+17, 1.288743972967732e+17, 1.288743973008358e+17, 1.288743973048982e+17, 1.288743973088045e+17, 1.288743973128669e+17, 1.288743973167732e+17, 1.288743973208358e+17, 1.288743973248982e+17, 1.288743973288045e+17, 1.288743973328669e+17, 1.288743973367732e+17, 1.288743973408357e+17, 1.288743973448983e+17, 1.288743973488046e+17, 1.288743973528669e+17, 1.288743973567732e+17, 1.288743973608357e+17, 1.288743973648982e+17, 1.288743973688045e+17, 1.288743973728669e+17, 1.288743973767732e+17, 1.288743973808357e+17, 1.288743973848983e+17, 1.288743973888045e+17, 1.288743973928671e+17, 1.288743973967732e+17, 1.288743974008357e+17, 1.288743974048983e+17, 1.288743974088045e+17, 1.288743974128669e+17, 1.288743974167732e+17, 1.288743974208357e+17, 1.288743974248983e+17, 1.288743974288045e+17, 1.288743974328671e+17, 1.288743974367732e+17, 1.288743974408357e+17, 1.288743974448983e+17, 1.288743974488045e+17, 1.288743974528671e+17, 1.288743974567732e+17, 1.288743974608357e+17, 1.288743974648983e+17, 1.288743974688045e+17, 1.288743974728671e+17, 1.288743974767732e+17, 1.288743974808357e+17, 1.288743974848983e+17, 1.288743974888045e+17, 1.288743974928671e+17, 1.288743974967732e+17, 1.288743975008357e+17, 1.288743975048983e+17, 1.288743975088045e+17, 1.288743975128671e+17, 1.288743975167732e+17, 1.288743975208358e+17, 1.288743975248983e+17, 1.288743975288045e+17, 1.288743975328671e+17, 1.288743975367732e+17, 1.288743975408357e+17, 1.288743975448982e+17, 1.288743975488045e+17, 1.288743975528671e+17, 1.288743975567732e+17, 1.288743975608358e+17, 1.288743975648982e+17, 1.288743975688045e+17, 1.288743975728669e+17, 1.288743975767732e+17, 1.288743975808358e+17, 1.288743975848982e+17, 1.288743975888045e+17, 1.288743975928669e+17, 1.288743975967732e+17, 1.288743976008357e+17, 1.288743976048983e+17, 1.288743976088046e+17, 1.288743976128669e+17, 1.288743976167732e+17, 1.288743976208357e+17, 1.288743976248982e+17, 1.288743976288045e+17, 1.288743976328669e+17, 1.288743976367732e+17, 1.288743976408357e+17, 1.288743976448983e+17, 1.288743976488045e+17, 1.288743976528671e+17, 1.288743976567732e+17, 1.288743976608357e+17, 1.288743976648983e+17, 1.288743976688045e+17, 1.288743976728669e+17, 1.288743976767732e+17, 1.288743976808357e+17, 1.288743976848983e+17, 1.288743976888045e+17, 1.288743976928671e+17, 1.288743976967732e+17, 1.288743977008357e+17, 1.288743977048983e+17, 1.288743977088045e+17, 1.288743977128671e+17, 1.288743977167731e+17, 1.288743977208357e+17, 1.288743977248983e+17, 1.288743977288045e+17, 1.288743977328671e+17, 1.288743977367732e+17, 1.288743977408357e+17, 1.288743977448983e+17, 1.288743977488045e+17, 1.288743977528671e+17, 1.288743977567732e+17, 1.288743977608357e+17, 1.288743977648983e+17, 1.288743977652407e+17, 1.288743977693033e+17, 1.288743977732095e+17, 1.288743977772719e+17, 1.288743977813345e+17, 1.288743977852407e+17, 1.288743977893033e+17, 1.288743977932095e+17, 1.288743977972721e+17, 1.288743978013345e+17, 1.288743978052407e+17, 1.288743978093033e+17, 1.288743978132095e+17, 1.288743978172719e+17, 1.288743978213345e+17, 1.288743978252407e+17, 1.288743978293033e+17, 1.288743978332095e+17, 1.288743978372721e+17, 1.288743978413345e+17, 1.288743978452408e+17, 1.288743978493033e+17, 1.288743978532095e+17, 1.288743978572721e+17, 1.288743978613344e+17, 1.288743978652407e+17, 1.288743978693033e+17, 1.288743978732095e+17, 1.288743978772721e+17, 1.288743978813345e+17, 1.288743978852408e+17, 1.288743978893032e+17, 1.288743978932095e+17, 1.288743978972721e+17, 1.288743979013344e+17, 1.288743979052408e+17, 1.288743979093032e+17, 1.288743979132095e+17, 1.288743979172719e+17, 1.288743979213345e+17, 1.288743979252408e+17, 1.288743979293032e+17, 1.288743979332096e+17, 1.288743979372719e+17, 1.288743979413345e+17, 1.288743979452407e+17, 1.288743979493032e+17, 1.288743979532095e+17, 1.288743979572719e+17, 1.288743979613345e+17, 1.288743979652407e+17, 1.288743979693033e+17, 1.288743979732095e+17, 1.288743979772719e+17, 1.288743979813345e+17, 1.288743979852407e+17, 1.288743979893032e+17, 1.288743979932095e+17, 1.288743979972719e+17, 1.288743980013345e+17, 1.288743980052407e+17, 1.288743980093033e+17, 1.288743980132095e+17, 1.288743980172721e+17, 1.288743980213345e+17, 1.288743980252407e+17, 1.288743980293033e+17, 1.288743980332095e+17, 1.288743980372719e+17, 1.288743980413345e+17, 1.288743980452407e+17, 1.288743980493033e+17, 1.288743980532095e+17, 1.288743980572721e+17, 1.288743980613345e+17, 1.288743980652407e+17, 1.288743980693033e+17, 1.288743980732095e+17, 1.288743980772721e+17, 1.288743980813345e+17, 1.288743980852407e+17, 1.288743980893033e+17, 1.288743980932095e+17, 1.288743980972721e+17, 1.288743981013344e+17, 1.288743981052408e+17, 1.288743981093033e+17, 1.288743981132095e+17, 1.288743981172721e+17, 1.288743981213344e+17, 1.288743981252407e+17, 1.288743981293032e+17, 1.288743981332095e+17, 1.288743981372721e+17, 1.288743981413345e+17, 1.288743981452408e+17, 1.288743981493032e+17, 1.288743981532095e+17, 1.288743981572719e+17, 1.288743981613344e+17, 1.288743981652408e+17, 1.288743981693032e+17, 1.288743981732095e+17, 1.288743981772719e+17, 1.288743981813345e+17, 1.288743981852407e+17, 1.288743981893032e+17, 1.288743981932096e+17, 1.288743981972719e+17, 1.288743982013345e+17, 1.288743982052407e+17, 1.288743982093032e+17, 1.288743982132095e+17, 1.288743982172719e+17, 1.288743982213345e+17, 1.288743982252407e+17, 1.288743982293033e+17, 1.288743982332095e+17, 1.288743982372719e+17, 1.288743982413345e+17, 1.288743982452407e+17, 1.288743982493032e+17, 1.288743982532095e+17, 1.288743982572719e+17, 1.288743982613345e+17, 1.288743982652407e+17, 1.288743982693033e+17, 1.288743982732095e+17, 1.288743982772721e+17, 1.288743982813345e+17, 1.288743982852407e+17, 1.288743982893033e+17, 1.288743982932095e+17, 1.288743982972719e+17, 1.288743983013345e+17, 1.288743983052407e+17, 1.288743983093033e+17, 1.288743983132095e+17, 1.288743983172721e+17, 1.288743983213345e+17, 1.288743983252407e+17, 1.288743983293033e+17, 1.288743983332095e+17, 1.288743983372721e+17, 1.288743983413345e+17, 1.288743983452407e+17, 1.288743983493033e+17, 1.288743983532095e+17, 1.288743983572721e+17, 1.288743983613344e+17, 1.288743983652408e+17, 1.288743983693033e+17, 1.288743983732095e+17, 1.288743983772721e+17, 1.288743983813344e+17, 1.288743983852407e+17, 1.288743983893032e+17, 1.288743983932095e+17, 1.288743983972721e+17, 1.288743984013345e+17, 1.288743984052408e+17, 1.288743984093032e+17, 1.288743984132096e+17, 1.288743984172719e+17, 1.288743984213344e+17, 1.288743984252408e+17, 1.288743984293032e+17, 1.288743984332095e+17, 1.288743984372719e+17, 1.288743984413345e+17, 1.288743984452407e+17, 1.288743984493033e+17, 1.288743984532096e+17, 1.288743984572719e+17, 1.288743984613345e+17, 1.288743984652407e+17, 1.288743984693032e+17, 1.288743984732095e+17, 1.288743984772719e+17, 1.288743984813345e+17, 1.288743984852407e+17, 1.288743984893033e+17, 1.288743984932095e+17, 1.288743984972719e+17, 1.288743985013345e+17, 1.288743985052407e+17, 1.288743985093033e+17, 1.288743985132095e+17, 1.288743985172719e+17, 1.288743985213345e+17, 1.288743985252407e+17, 1.288743985293033e+17, 1.288743985332095e+17, 1.288743985372721e+17, 1.288743985413345e+17, 1.288743985452407e+17, 1.288743985493033e+17, 1.288743985532095e+17, 1.288743985572719e+17, 1.288743985613345e+17, 1.288743985652407e+17, 1.288743985693033e+17, 1.288743985732095e+17, 1.288743985772721e+17, 1.288743985813345e+17, 1.288743985852407e+17, 1.288743985893033e+17, 1.288743985932095e+17, 1.288743985972721e+17, 1.288743986013345e+17, 1.288743986052407e+17, 1.288743986093033e+17, 1.288743986132095e+17, 1.288743986172721e+17, 1.288743986213344e+17, 1.288743986252408e+17, 1.288743986293033e+17, 1.288743986332095e+17, 1.288743986372721e+17, 1.288743986413344e+17, 1.288743986452407e+17, 1.288743986493032e+17, 1.288743986532095e+17, 1.288743986572721e+17, 1.288743986613345e+17, 1.288743986652408e+17, 1.288743986693032e+17, 1.288743986732096e+17, 1.288743986772719e+17, 1.288743986813344e+17, 1.288743986852408e+17, 1.288743986893032e+17, 1.288743986932095e+17, 1.288743986972719e+17, 1.288743987013345e+17, 1.288743987052407e+17, 1.288743987093033e+17, 1.288743987132096e+17, 1.288743987172719e+17, 1.288743987213345e+17, 1.288743987252407e+17, 1.288743987293032e+17, 1.288743987332095e+17, 1.288743987372719e+17, 1.288743987413345e+17, 1.288743987452407e+17, 1.288743987493033e+17, 1.288743987532095e+17, 1.288743987572719e+17, 1.288743987613345e+17, 1.288743987652407e+17, 1.288743987693033e+17, 1.288743987732095e+17, 1.288743987772719e+17, 1.288743987813345e+17, 1.288743987852407e+17, 1.288743987893033e+17, 1.288743987932095e+17, 1.288743987972721e+17, 1.288743988013345e+17, 1.288743988052407e+17, 1.288743988093033e+17, 1.288743988132095e+17, 1.288743988172719e+17, 1.288743988213345e+17, 1.288743988252407e+17, 1.288743988293033e+17, 1.288743988332095e+17, 1.288743988372721e+17, 1.288743988413345e+17, 1.288743988452407e+17, 1.288743988493033e+17, 1.288743988532095e+17, 1.288743988572721e+17, 1.288743988613345e+17, 1.288743988652407e+17, 1.288743988693033e+17, 1.288743988732095e+17, 1.288743988772721e+17, 1.288743988813345e+17, 1.288743988852408e+17, 1.288743988893033e+17, 1.288743988932095e+17, 1.288743988972721e+17, 1.288743989013344e+17, 1.288743989052407e+17, 1.288743989093032e+17, 1.288743989132095e+17, 1.288743989172721e+17, 1.288743989213345e+17, 1.288743989252408e+17, 1.288743989293032e+17, 1.288743989332096e+17, 1.288743989372719e+17, 1.288743989413344e+17, 1.288743989452408e+17, 1.288743989493032e+17, 1.288743989532095e+17, 1.288743989572719e+17, 1.288743989613345e+17, 1.288743989652407e+17, 1.288743989693033e+17, 1.288743989732096e+17, 1.288743989772719e+17, 1.288743989813345e+17, 1.288743989852407e+17, 1.288743989893032e+17, 1.288743989932095e+17, 1.288743989972719e+17, 1.288743990013345e+17, 1.288743990052407e+17, 1.288743990093033e+17, 1.288743990132095e+17, 1.288743990172719e+17, 1.288743990213345e+17, 1.288743990252407e+17, 1.288743990293033e+17, 1.288743990332095e+17, 1.288743990372719e+17, 1.288743990413345e+17, 1.288743990452407e+17, 1.288743990493033e+17, 1.288743990532095e+17, 1.288743990572721e+17, 1.288743990613345e+17, 1.288743990652407e+17, 1.288743990693033e+17, 1.288743990732095e+17, 1.288743990772719e+17, 1.288743990813345e+17, 1.288743990852407e+17, 1.288743990893033e+17, 1.288743990932095e+17, 1.288743990972721e+17, 1.288743991013345e+17, 1.288743991052408e+17, 1.288743991093033e+17, 1.288743991132095e+17, 1.288743991172721e+17, 1.288743991213344e+17, 1.288743991252407e+17, 1.288743991293033e+17, 1.288743991332095e+17, 1.288743991372721e+17, 1.288743991413345e+17, 1.288743991452408e+17, 1.288743991493032e+17, 1.288743991532095e+17, 1.288743991572721e+17, 1.288743991613344e+17, 1.288743991652408e+17, 1.288743991693032e+17, 1.288743991732095e+17, 1.288743991772719e+17, 1.288743991813345e+17, 1.288743991852408e+17, 1.288743991893032e+17, 1.288743991932096e+17, 1.288743991972719e+17, 1.288743992013345e+17, 1.288743992052407e+17, 1.288743992093032e+17, 1.288743992132095e+17, 1.288743992172719e+17, 1.288743992213345e+17, 1.288743992252407e+17, 1.288743992293033e+17, 1.288743992332095e+17, 1.288743992372719e+17, 1.288743992413345e+17, 1.288743992452407e+17, 1.288743992493032e+17, 1.288743992532095e+17, 1.288743992572719e+17, 1.288743992613345e+17, 1.288743992652407e+17, 1.288743992693033e+17, 1.288743992732095e+17, 1.288743992772719e+17, 1.288743992813345e+17, 1.288743992932095e+17, 1.288743992972719e+17, 1.288743993013345e+17, 1.288743993052407e+17, 1.288743993093033e+17, 1.288743993132095e+17, 1.288743993172721e+17, 1.288743993213345e+17, 1.288743993252407e+17, 1.288743993293033e+17, 1.288743993332095e+17, 1.288743993372719e+17, 1.288743993413345e+17, 1.288743993452407e+17, 1.288743993493033e+17, 1.288743993532095e+17, 1.288743993572721e+17, 1.288743993613345e+17, 1.288743993652408e+17, 1.288743993693033e+17, 1.288743993732095e+17, 1.288743993772721e+17, 1.288743993813344e+17, 1.288743993852407e+17, 1.288743993893033e+17, 1.288743993932095e+17, 1.288743993972721e+17, 1.288743994013345e+17, 1.288743994052408e+17, 1.288743994093032e+17, 1.288743994132095e+17, 1.288743994172721e+17, 1.288743994213344e+17, 1.288743994252408e+17, 1.288743994293032e+17, 1.288743994332095e+17, 1.288743994372719e+17, 1.288743994413345e+17, 1.288743994452408e+17, 1.288743994493032e+17, 1.288743994532096e+17, 1.288743994572719e+17, 1.288743994613345e+17, 1.288743994652407e+17, 1.288743994693032e+17, 1.288743994732095e+17, 1.288743994772719e+17, 1.288743994813345e+17, 1.288743994852407e+17, 1.288743994893033e+17, 1.288743994932095e+17, 1.288743994972719e+17, 1.288743995013345e+17, 1.288743995052407e+17, 1.288743995093032e+17, 1.288743995132095e+17, 1.288743995172719e+17, 1.288743995213345e+17, 1.288743995252407e+17, 1.288743995293033e+17, 1.288743995332095e+17, 1.288743995372719e+17, 1.288743995413345e+17, 1.288743995452407e+17, 1.288743995493033e+17, 1.288743995532095e+17, 1.288743995572719e+17, 1.288743995613345e+17, 1.288743995652407e+17, 1.288743995693033e+17, 1.288743995732095e+17, 1.288743995772721e+17, 1.288743995813345e+17, 1.288743995852407e+17, 1.288743995893033e+17, 1.288743995932095e+17, 1.288743995972719e+17, 1.288743996013345e+17, 1.288743996052407e+17, 1.288743996093033e+17, 1.288743996132095e+17, 1.288743996172721e+17, 1.288743996213345e+17, 1.288743996252408e+17, 1.288743996293033e+17, 1.288743996332095e+17, 1.288743996372721e+17, 1.288743996413344e+17, 1.288743996452407e+17, 1.288743996493033e+17, 1.288743996532095e+17, 1.288743996572721e+17, 1.288743996613345e+17, 1.288743996652408e+17, 1.288743996693032e+17, 1.288743996732095e+17, 1.288743996772721e+17, 1.288743996813344e+17, 1.288743996852408e+17, 1.288743996893032e+17, 1.288743996932095e+17, 1.288743996972719e+17, 1.288743997013345e+17, 1.288743997052408e+17, 1.288743997093032e+17, 1.288743997132096e+17, 1.288743997172719e+17, 1.288743997213345e+17, 1.288743997252407e+17, 1.288743997293032e+17, 1.288743997332095e+17, 1.288743997372719e+17, 1.288743997413345e+17, 1.288743997452407e+17, 1.288743997493033e+17, 1.288743997532095e+17, 1.288743997572719e+17, 1.288743997613345e+17, 1.288743997652407e+17, 1.288743997693032e+17, 1.288743997732095e+17, 1.288743997772719e+17, 1.288743997813345e+17, 1.288743997852407e+17, 1.288743997893033e+17, 1.288743997932095e+17, 1.288743997972721e+17, 1.288743998013345e+17, 1.288743998052407e+17, 1.288743998093033e+17, 1.288743998132095e+17, 1.288743998172719e+17, 1.288743998213345e+17, 1.288743998252407e+17, 1.288743998293033e+17, 1.288743998332095e+17, 1.288743998372721e+17, 1.288743998413345e+17, 1.288743998452407e+17, 1.288743998493033e+17, 1.288743998532095e+17, 1.288743998572721e+17, 1.288743998613345e+17, 1.288743998652407e+17, 1.288743998693033e+17, 1.288743998732095e+17, 1.288743998772721e+17, 1.288743998813345e+17, 1.288743998852408e+17, 1.288743998893033e+17, 1.288743998932095e+17, 1.288743998972721e+17, 1.288743999013344e+17, 1.288743999052407e+17, 1.288743999093033e+17, 1.288743999132095e+17, 1.288743999172721e+17, 1.288743999213345e+17, 1.288743999252408e+17, 1.288743999293032e+17, 1.288743999332095e+17, 1.288743999372721e+17, 1.288743999413344e+17, 1.288743999452408e+17, 1.288743999493032e+17, 1.288743999532095e+17, 1.288743999572719e+17, 1.288743999613345e+17, 1.288743999652408e+17, 1.288743999693032e+17, 1.288743999732096e+17, 1.288743999772719e+17, 1.288743999813345e+17, 1.288743999852407e+17, 1.288743999893032e+17, 1.288743999932095e+17, 1.288743999972719e+17, 1.288744000013345e+17, 1.288744000052407e+17, 1.288744000172719e+17, 1.288744000213345e+17, 1.288744000252407e+17, 1.288744000293032e+17, 1.288744000332095e+17, 1.288744000372719e+17, 1.288744000413345e+17, 1.288744000452407e+17, 1.288744000493033e+17, 1.288744000532095e+17, 1.288744000572721e+17, 1.288744000613345e+17, 1.288744000652407e+17, 1.288744000693033e+17, 1.288744000732095e+17, 1.288744000813345e+17, 1.288744000852407e+17, 1.288744000893033e+17, 1.288744000932095e+17, 1.288744000972721e+17, 1.288744001013345e+17, 1.288744001052407e+17, 1.288744001093033e+17, 1.288744001132095e+17, 1.288744001213345e+17, 1.288744001252407e+17, 1.288744001293033e+17, 1.288744001332095e+17, 1.288744001372721e+17, 1.288744001413344e+17, 1.288744001452408e+17, 1.288744001493033e+17, 1.288744001532095e+17, 1.288744001572721e+17, 1.288744001613344e+17, 1.288744001652407e+17, 1.288744001693032e+17, 1.288744001732095e+17, 1.288744001772721e+17, 1.288744001813345e+17, 1.288744001852408e+17, 1.288744001893032e+17, 1.288744002093032e+17, 1.288744002213345e+17, 1.288744002252407e+17, 1.288744002293033e+17, 1.288744002332096e+17, 1.288744002372719e+17, 1.288744002413345e+17, 1.288744002452407e+17, 1.288744002493032e+17, 1.288744002532095e+17, 1.288744002572719e+17, 1.288744002613345e+17, 1.288744002652407e+17, 1.288744002693033e+17, 1.288744002732095e+17, 1.288744002772719e+17, 1.288744002813345e+17, 1.288744002852407e+17, 1.288744002893032e+17, 1.288744002932095e+17, 1.288744002972719e+17, 1.288744003013345e+17, 1.288744003052407e+17, 1.288744003093033e+17, 1.288744003132095e+17, 1.288744003172721e+17, 1.288744003213345e+17, 1.288744003252407e+17, 1.288744003293033e+17, 1.288744003332095e+17, 1.288744003372719e+17, 1.288744003413345e+17, 1.288744003452407e+17, 1.288744003532095e+17, 1.288744003572721e+17, 1.288744003613345e+17, 1.288744003652407e+17, 1.288744003693033e+17, 1.288744003732095e+17, 1.288744003772721e+17, 1.288744003813345e+17, 1.288744003852407e+17, 1.288744003893033e+17, 1.288744003932095e+17, 1.288744003972721e+17, 1.288744004013344e+17, 1.288744004052408e+17, 1.288744004093033e+17, 1.288744004132095e+17, 1.288744004172721e+17, 1.288744004213344e+17, 1.288744004252407e+17, 1.288744004293032e+17, 1.288744004332095e+17, 1.288744004452408e+17, 1.288744004532096e+17, 1.288744004572719e+17, 1.288744004613344e+17, 1.288744004652408e+17, 1.288744004693032e+17, 1.288744004732095e+17, 1.288744004772719e+17, 1.288744004852407e+17, 1.288744004893033e+17, 1.288744004932096e+17, 1.288744004972719e+17, 1.288744005013345e+17, 1.288744005052407e+17, 1.288744005093032e+17, 1.288744005132095e+17, 1.288744005172719e+17, 1.288744005213345e+17, 1.288744005252407e+17, 1.288744005293033e+17, 1.288744005332095e+17, 1.288744005372719e+17, 1.288744005413345e+17, 1.288744005452407e+17, 1.288744005493033e+17, 1.288744005532095e+17, 1.288744005572719e+17, 1.288744005613345e+17, 1.288744005652407e+17, 1.288744005693033e+17, 1.288744005732095e+17, 1.288744005772721e+17, 1.288744005813345e+17, 1.288744005852407e+17, 1.288744005893033e+17, 1.288744005932095e+17, 1.288744005972719e+17, 1.288744006013345e+17, 1.288744006052407e+17, 1.288744006093033e+17, 1.288744006132095e+17, 1.288744006172721e+17, 1.288744006213345e+17, 1.288744006252407e+17, 1.288744006293033e+17, 1.288744006372721e+17, 1.288744006413345e+17, 1.288744006452407e+17, 1.288744006493033e+17, 1.288744006532095e+17, 1.288744006572721e+17, 1.288744006613344e+17, 1.288744006652408e+17, 1.288744006693033e+17, 1.288744006732095e+17, 1.288744006772721e+17, 1.288744006813344e+17, 1.288744006852407e+17, 1.288744006893032e+17, 1.288744006932095e+17, 1.288744006972721e+17, 1.288744007013345e+17, 1.288744007052408e+17, 1.288744007093032e+17, 1.288744007132096e+17, 1.288744007252408e+17, 1.288744007293032e+17, 1.288744007332095e+17, 1.288744007372719e+17, 1.288744007413345e+17, 1.288744007452407e+17, 1.288744007493033e+17, 1.288744007532096e+17, 1.288744007572719e+17, 1.288744007613345e+17, 1.288744007652407e+17, 1.288744007693032e+17, 1.288744007732095e+17, 1.288744007772719e+17, 1.288744007813345e+17, 1.288744007852407e+17, 1.288744007893033e+17, 1.288744007932095e+17, 1.288744007972719e+17, 1.288744008013345e+17, 1.288744008052407e+17, 1.288744008093033e+17, 1.288744008132095e+17, 1.288744008172719e+17, 1.288744008213345e+17, 1.288744008252407e+17, 1.288744008293033e+17, 1.288744008332095e+17, 1.288744008372721e+17, 1.288744008413345e+17, 1.288744008452407e+17, 1.288744008493033e+17, 1.288744008532095e+17, 1.288744008572719e+17, 1.288744008613345e+17, 1.288744008652407e+17, 1.288744008693033e+17, 1.288744008732095e+17, 1.288744008772721e+17, 1.288744008813345e+17, 1.288744008852408e+17, 1.288744008893033e+17, 1.288744008932095e+17, 1.288744008972721e+17, 1.288744009013345e+17, 1.288744009052407e+17, 1.288744009093033e+17, 1.288744009132095e+17, 1.288744009172721e+17, 1.288744009213345e+17, 1.288744009252408e+17, 1.288744009293033e+17, 1.288744009332095e+17, 1.288744009372721e+17, 1.288744009413344e+17, 1.288744009452407e+17, 1.288744009493032e+17, 1.288744009532095e+17, 1.288744009572721e+17, 1.288744009613345e+17, 1.288744009652408e+17, 1.288744009693032e+17, 1.288744009732096e+17, 1.288744009772719e+17, 1.288744009813344e+17, 1.288744009852408e+17, 1.288744009893032e+17, 1.288744009932095e+17, 1.288744009972719e+17, 1.288744010013345e+17, 1.288744010052407e+17, 1.288744010093033e+17, 1.288744010132096e+17, 1.288744010172719e+17, 1.288744010213345e+17, 1.288744010252407e+17, 1.288744010293032e+17, 1.288744010332095e+17, 1.288744010372719e+17, 1.288744010413345e+17, 1.288744010452407e+17, 1.288744010493033e+17, 1.288744010532095e+17, 1.288744010572719e+17, 1.288744010613345e+17, 1.288744010652407e+17, 1.288744010693033e+17, 1.288744010732095e+17, 1.288744010772719e+17, 1.288744010813345e+17, 1.288744010852407e+17, 1.288744010893033e+17, 1.288744010932095e+17, 1.288744010972721e+17, 1.288744011013345e+17, 1.288744011052407e+17, 1.288744011093033e+17, 1.288744011132095e+17, 1.288744011172719e+17, 1.288744011213345e+17, 1.288744011252407e+17, 1.288744011293033e+17, 1.288744011332095e+17, 1.288744011372721e+17, 1.288744011413345e+17, 1.288744011452408e+17, 1.288744011493033e+17, 1.288744011532095e+17, 1.288744011572721e+17, 1.288744011613344e+17, 1.288744011652407e+17, 1.288744011693033e+17, 1.288744011732095e+17, 1.288744011772721e+17, 1.288744011813345e+17, 1.288744011852408e+17, 1.288744011893032e+17, 1.288744011932095e+17, 1.288744011972721e+17, 1.288744012013344e+17, 1.288744012052408e+17, 1.288744012093032e+17, 1.288744012132095e+17, 1.288744012172719e+17, 1.288744012213345e+17, 1.288744012252408e+17, 1.288744012293032e+17, 1.288744012332096e+17, 1.288744012372719e+17, 1.288744012413345e+17, 1.288744012452407e+17, 1.288744012493032e+17, 1.288744012532095e+17, 1.288744012572719e+17, 1.288744012613345e+17, 1.288744012652407e+17, 1.288744012693033e+17, 1.288744012732095e+17, 1.288744012772719e+17, 1.288744012813345e+17, 1.288744012852407e+17, 1.288744012893032e+17, 1.288744012932095e+17, 1.288744012972719e+17, 1.288744013013345e+17, 1.288744013052407e+17, 1.288744013093033e+17, 1.288744013132095e+17, 1.288744013172719e+17, 1.288744013213345e+17, 1.288744013252407e+17, 1.288744013293033e+17, 1.288744013332095e+17, 1.288744013372719e+17, 1.288744013413345e+17, 1.288744013452407e+17, 1.288744013493033e+17, 1.288744013532095e+17, 1.288744013572721e+17, 1.288744013613345e+17, 1.288744013652407e+17, 1.288744013693033e+17, 1.288744013732095e+17, 1.288744013772719e+17, 1.288744013813345e+17, 1.288744013852407e+17, 1.288744013893033e+17, 1.288744013932095e+17, 1.288744013972721e+17, 1.288744014013345e+17, 1.288744014052408e+17, 1.288744014093033e+17, 1.288744014132095e+17, 1.288744014172721e+17, 1.288744014213344e+17, 1.288744014252407e+17, 1.288744014293033e+17, 1.288744014332095e+17, 1.288744014372721e+17, 1.288744014413345e+17, 1.288744014452408e+17, 1.288744014493032e+17, 1.288744014532095e+17, 1.288744014572721e+17, 1.288744014613344e+17, 1.288744014652408e+17, 1.288744014693032e+17, 1.288744014732095e+17, 1.288744014772719e+17, 1.288744014813345e+17, 1.288744014852408e+17, 1.288744014893032e+17, 1.288744014932096e+17, 1.288744014972719e+17, 1.288744015013345e+17, 1.288744015052407e+17, 1.288744015093032e+17, 1.288744015132095e+17, 1.288744015172719e+17, 1.288744015213345e+17, 1.288744015252407e+17, 1.288744015293033e+17, 1.288744015332095e+17, 1.288744015372719e+17, 1.288744015413345e+17, 1.288744015452407e+17, 1.288744015493032e+17, 1.288744015532095e+17, 1.288744015572719e+17, 1.288744015613345e+17, 1.288744015652407e+17, 1.288744015693033e+17, 1.288744015732095e+17, 1.288744015772721e+17, 1.288744015813345e+17, 1.288744015852407e+17, 1.288744015893033e+17, 1.288744015932095e+17, 1.288744015972719e+17, 1.288744016013345e+17, 1.288744016052407e+17, 1.288744016093033e+17, 1.288744016132095e+17, 1.288744016172721e+17, 1.288744016213345e+17, 1.288744016252407e+17, 1.288744016293033e+17, 1.288744016332095e+17, 1.288744016372719e+17, 1.288744016413345e+17, 1.288744016452407e+17, 1.288744016493033e+17, 1.288744016532095e+17, 1.288744016572721e+17, 1.288744016613345e+17, 1.288744016652408e+17, 1.288744016693033e+17, 1.288744016732095e+17, 1.288744016772721e+17, 1.288744016813344e+17, 1.288744016852407e+17, 1.288744016893033e+17, 1.288744016932095e+17, 1.288744016972721e+17, 1.288744017013345e+17, 1.288744017052408e+17, 1.288744017093032e+17, 1.288744017132095e+17, 1.288744017172721e+17, 1.288744017213344e+17, 1.288744017252408e+17, 1.288744017293032e+17, 1.288744017332095e+17, 1.288744017372719e+17, 1.288744017413345e+17, 1.288744017452408e+17, 1.288744017493032e+17, 1.288744017532096e+17, 1.288744017572719e+17, 1.288744017613345e+17, 1.288744017652407e+17, 1.288744017693032e+17, 1.288744017732095e+17, 1.288744017772719e+17, 1.288744017813345e+17, 1.288744017852407e+17, 1.288744017893033e+17, 1.288744017932095e+17, 1.288744017972719e+17, 1.288744018013345e+17, 1.288744018052407e+17, 1.288744018093032e+17, 1.288744018132095e+17, 1.288744018172719e+17, 1.288744018213345e+17, 1.288744018252407e+17, 1.288744018293033e+17, 1.288744018332095e+17, 1.288744018372721e+17, 1.288744018413345e+17, 1.288744018452407e+17, 1.288744018493033e+17, 1.288744018532095e+17, 1.288744018572719e+17, 1.288744018613345e+17, 1.288744018652407e+17, 1.288744018693033e+17, 1.288744018732095e+17, 1.288744018772721e+17, 1.288744018813345e+17, 1.288744018852407e+17, 1.288744018893033e+17, 1.288744018932095e+17, 1.288744018972721e+17, 1.288744019013345e+17, 1.288744019052407e+17, 1.288744019093033e+17, 1.288744019132095e+17, 1.288744019172721e+17, 1.288744019213345e+17, 1.288744019252408e+17, 1.288744019293033e+17, 1.288744019332095e+17, 1.288744019372721e+17, 1.288744019413344e+17, 1.288744019452407e+17, 1.288744019493033e+17, 1.288744019532095e+17, 1.288744019572721e+17, 1.288744019613345e+17, 1.288744019652408e+17, 1.288744019693032e+17, 1.288744019732095e+17, 1.288744019772721e+17, 1.288744019813344e+17, 1.288744019852408e+17, 1.288744019893032e+17, 1.288744019932095e+17, 1.288744019972719e+17, 1.288744020013345e+17, 1.288744020052408e+17, 1.288744020093032e+17, 1.288744020132096e+17, 1.288744020172719e+17, 1.288744020213345e+17, 1.288744020252407e+17, 1.288744020293032e+17, 1.288744020332095e+17, 1.288744020372719e+17, 1.288744020413345e+17, 1.288744020452407e+17, 1.288744020493033e+17, 1.288744020532095e+17, 1.288744020572719e+17, 1.288744020613345e+17, 1.288744020652407e+17, 1.288744020693032e+17, 1.288744020732095e+17, 1.288744020772719e+17, 1.288744020813345e+17, 1.288744020852407e+17, 1.288744020893033e+17, 1.288744020932095e+17, 1.288744020972721e+17, 1.288744021013345e+17, 1.288744021052407e+17, 1.288744021093033e+17, 1.288744021132095e+17, 1.288744021172719e+17, 1.288744021213345e+17, 1.288744021252407e+17, 1.288744021293033e+17, 1.288744021332095e+17, 1.288744021372721e+17, 1.288744021413345e+17, 1.288744021452407e+17, 1.288744021493033e+17, 1.288744021532095e+17, 1.288744021572721e+17, 1.288744021613345e+17, 1.288744021652407e+17, 1.288744021693033e+17, 1.288744021732095e+17, 1.288744021772721e+17, 1.288744021813344e+17, 1.288744021852408e+17, 1.288744021893033e+17, 1.288744021932095e+17, 1.288744021972721e+17, 1.288744022013344e+17, 1.288744022052407e+17, 1.288744022093032e+17, 1.288744022132095e+17, 1.288744022172721e+17, 1.288744022213345e+17, 1.288744022252408e+17, 1.288744022293032e+17, 1.288744022332096e+17, 1.288744022372719e+17, 1.288744022413344e+17, 1.288744022452408e+17, 1.288744022493032e+17, 1.288744022532095e+17, 1.288744022572719e+17, 1.288744022613345e+17, 1.288744022652407e+17, 1.288744022693033e+17, 1.288744022732096e+17, 1.288744022772719e+17, 1.288744022813345e+17, 1.288744022852407e+17, 1.288744022893032e+17, 1.288744022932095e+17, 1.288744022972719e+17, 1.288744023013345e+17, 1.288744023052407e+17, 1.288744023093033e+17, 1.288744023132095e+17, 1.288744023172719e+17, 1.288744023213345e+17, 1.288744023252407e+17, 1.288744023293033e+17, 1.288744023332095e+17, 1.288744023372719e+17, 1.288744023413345e+17, 1.288744023452407e+17, 1.288744023493033e+17, 1.288744023532095e+17, 1.288744023572721e+17, 1.288744023613345e+17, 1.288744023652407e+17, 1.288744023693033e+17, 1.288744023732095e+17, 1.288744023772719e+17, 1.288744023813345e+17, 1.288744023852407e+17, 1.288744023893033e+17, 1.288744023932095e+17, 1.288744023972721e+17, 1.288744024013345e+17, 1.288744024052407e+17, 1.288744024093033e+17, 1.288744024132095e+17, 1.288744024172721e+17, 1.288744024213345e+17, 1.288744024252407e+17, 1.288744024293033e+17, 1.288744024332095e+17, 1.288744024372721e+17, 1.288744024413344e+17, 1.288744024452408e+17, 1.288744024493033e+17, 1.288744024532095e+17, 1.288744024572721e+17, 1.288744024613344e+17, 1.288744024652407e+17, 1.288744024693032e+17, 1.288744024732095e+17, 1.288744024772721e+17, 1.288744024813345e+17, 1.288744024852408e+17, 1.288744024893032e+17, 1.288744024932096e+17, 1.288744024972719e+17, 1.288744025013344e+17, 1.288744025052408e+17, 1.288744025093032e+17, 1.288744025132095e+17, 1.288744025172719e+17, 1.288744025213345e+17, 1.288744025252407e+17, 1.288744025293033e+17, 1.288744025332096e+17, 1.288744025372719e+17, 1.288744025413345e+17, 1.288744025452407e+17, 1.288744025493032e+17, 1.288744025532095e+17, 1.288744025572719e+17, 1.288744025613345e+17, 1.288744025652407e+17, 1.288744025693033e+17, 1.288744025732095e+17, 1.288744025772719e+17, 1.288744025813345e+17, 1.288744025852407e+17, 1.288744025893033e+17, 1.288744025932095e+17, 1.288744025972719e+17, 1.288744026013345e+17, 1.288744026052407e+17, 1.288744026093033e+17, 1.288744026132095e+17, 1.288744026172721e+17, 1.288744026213345e+17, 1.288744026252407e+17, 1.288744026293033e+17, 1.288744026332095e+17, 1.288744026372719e+17, 1.288744026413345e+17, 1.288744026452407e+17, 1.288744026493033e+17, 1.288744026532095e+17, 1.288744026572721e+17, 1.288744026613345e+17, 1.288744026652407e+17, 1.288744026693033e+17, 1.288744026732095e+17, 1.288744026772721e+17, 1.288744026813345e+17, 1.288744026852407e+17, 1.288744026893033e+17, 1.288744026932095e+17, 1.288744026972721e+17, 1.288744027013344e+17, 1.288744027052408e+17, 1.288744027093033e+17, 1.288744027132095e+17, 1.288744027172721e+17, 1.288744027213344e+17, 1.288744027252407e+17, 1.288744027293032e+17, 1.288744027332095e+17, 1.288744027372721e+17, 1.288744027413345e+17, 1.288744027452408e+17, 1.288744027493032e+17, 1.288744027532096e+17, 1.288744027572719e+17, 1.288744027613344e+17, 1.288744027652408e+17, 1.288744027693032e+17, 1.288744027732095e+17, 1.288744027772719e+17, 1.288744027813345e+17, 1.288744027852407e+17, 1.288744027893033e+17, 1.288744027932096e+17, 1.288744027972719e+17, 1.288744028013345e+17, 1.288744028052407e+17, 1.288744028093032e+17, 1.288744028132095e+17, 1.288744028172719e+17, 1.288744028213345e+17, 1.288744028252407e+17, 1.288744028293033e+17, 1.288744028332095e+17, 1.288744028372719e+17, 1.288744028413345e+17, 1.288744028452407e+17, 1.288744028493033e+17, 1.288744028532095e+17, 1.288744028572719e+17, 1.288744028613345e+17, 1.288744028652407e+17, 1.288744028693033e+17, 1.288744028732095e+17, 1.288744028772721e+17, 1.288744028813345e+17, 1.288744028852407e+17, 1.288744028893033e+17, 1.288744028932095e+17, 1.288744028972719e+17, 1.288744029013345e+17, 1.288744029052407e+17, 1.288744029093033e+17, 1.288744029132095e+17, 1.288744029172721e+17, 1.288744029213345e+17, 1.288744029252408e+17, 1.288744029293033e+17, 1.288744029332095e+17, 1.288744029372721e+17, 1.288744029413344e+17, 1.288744029452407e+17, 1.288744029493033e+17, 1.288744029532095e+17, 1.288744029572721e+17, 1.288744029613345e+17, 1.288744029652408e+17, 1.288744029693032e+17, 1.288744029732095e+17, 1.288744029772721e+17, 1.288744029813344e+17, 1.288744029852407e+17, 1.288744029893032e+17, 1.288744029932095e+17, 1.288744029972719e+17, 1.288744030013345e+17, 1.288744030052408e+17, 1.288744030093032e+17, 1.288744030132096e+17, 1.288744030172719e+17, 1.288744030213345e+17, 1.288744030252407e+17, 1.288744030293032e+17, 1.288744030332095e+17, 1.288744030372719e+17, 1.288744030413345e+17, 1.288744030452407e+17, 1.288744030493033e+17, 1.288744030532095e+17, 1.288744030572719e+17, 1.288744030613345e+17, 1.288744030652407e+17, 1.288744030693032e+17, 1.288744030732095e+17, 1.288744030772719e+17, 1.288744030813345e+17, 1.288744030852407e+17, 1.288744030893033e+17, 1.288744030932095e+17, 1.288744030972719e+17, 1.288744031013345e+17, 1.288744031052407e+17, 1.288744031093033e+17, 1.288744031132095e+17, 1.288744031172719e+17, 1.288744031213345e+17, 1.288744031252407e+17, 1.288744031293033e+17, 1.288744031332095e+17, 1.288744031372721e+17, 1.288744031413345e+17, 1.288744031452407e+17, 1.288744031493033e+17, 1.288744031532095e+17, 1.288744031572719e+17, 1.288744031613345e+17, 1.288744031652407e+17, 1.288744031693033e+17, 1.288744031732095e+17, 1.288744031772721e+17, 1.288744031813345e+17, 1.288744031852408e+17, 1.288744031893033e+17, 1.288744031932095e+17, 1.288744031972721e+17, 1.288744032013344e+17, 1.288744032052407e+17, 1.288744032093033e+17, 1.288744032132095e+17, 1.288744032172721e+17, 1.288744032213345e+17, 1.288744032252408e+17, 1.288744032293032e+17, 1.288744032332095e+17, 1.288744032372721e+17, 1.288744032413344e+17, 1.288744032452408e+17, 1.288744032493032e+17, 1.288744032532095e+17, 1.288744032572719e+17, 1.288744032613345e+17, 1.288744032652408e+17, 1.288744032693032e+17, 1.288744032732096e+17, 1.288744032772719e+17, 1.288744032813345e+17, 1.288744032852407e+17, 1.288744032893032e+17, 1.288744032932095e+17, 1.288744032972719e+17, 1.288744033013345e+17, 1.288744033052407e+17, 1.288744033093033e+17, 1.288744033132095e+17, 1.288744033172719e+17, 1.288744033213345e+17, 1.288744033252407e+17, 1.288744033293032e+17, 1.288744033332095e+17, 1.288744033372719e+17, 1.288744033413345e+17, 1.288744033452407e+17, 1.288744033493033e+17, 1.288744033532095e+17, 1.288744033572719e+17, 1.288744033613345e+17, 1.288744033652407e+17, 1.288744033693033e+17, 1.288744033732095e+17, 1.288744033772719e+17, 1.288744033813345e+17, 1.288744033852407e+17, 1.288744033893033e+17, 1.288744033932095e+17, 1.288744033972721e+17, 1.288744034013345e+17, 1.288744034052407e+17, 1.288744034093033e+17, 1.288744034132095e+17, 1.288744034172719e+17, 1.288744034213345e+17, 1.288744034252407e+17, 1.288744034293033e+17, 1.288744034332095e+17, 1.288744034372721e+17, 1.288744034413345e+17, 1.288744034452408e+17, 1.288744034493033e+17, 1.288744034532095e+17, 1.288744034572721e+17, 1.288744034613344e+17, 1.288744034652407e+17, 1.288744034693033e+17, 1.288744034732095e+17, 1.288744034772721e+17, 1.288744034813345e+17, 1.288744034852408e+17, 1.288744034893032e+17, 1.288744034932095e+17, 1.288744034972721e+17, 1.288744035013344e+17, 1.288744035052408e+17, 1.288744035093032e+17, 1.288744035132095e+17, 1.288744035172719e+17, 1.288744035213345e+17, 1.288744035252408e+17, 1.288744035293032e+17, 1.288744035332096e+17, 1.288744035372719e+17, 1.288744035413345e+17, 1.288744035452407e+17, 1.288744035493032e+17, 1.288744035532095e+17, 1.288744035572719e+17, 1.288744035613345e+17, 1.288744035652407e+17, 1.288744035693033e+17, 1.288744035732095e+17, 1.288744035772719e+17, 1.288744035813345e+17, 1.288744035852407e+17, 1.288744035893032e+17, 1.288744035932095e+17, 1.288744035972719e+17, 1.288744036013345e+17, 1.288744036052407e+17, 1.288744036093033e+17, 1.288744036132095e+17, 1.288744036172721e+17, 1.288744036213345e+17, 1.288744036252407e+17, 1.288744036293033e+17, 1.288744036332095e+17, 1.288744036372719e+17, 1.288744036413345e+17, 1.288744036452407e+17, 1.288744036493033e+17, 1.288744036532095e+17, 1.288744036572721e+17, 1.288744036613345e+17, 1.288744036652407e+17, 1.288744036693033e+17, 1.288744036732095e+17, 1.288744036772721e+17, 1.288744036813345e+17, 1.288744036852407e+17, 1.288744036893033e+17, 1.288744036932095e+17, 1.288744036972721e+17, 1.288744037013345e+17, 1.288744037052408e+17, 1.288744037093033e+17, 1.288744037132095e+17, 1.288744037172721e+17, 1.288744037213344e+17, 1.288744037252407e+17, 1.288744037293033e+17, 1.288744037332095e+17, 1.288744037372721e+17, 1.288744037413345e+17, 1.288744037452408e+17, 1.288744037493032e+17, 1.288744037532095e+17, 1.288744037572721e+17, 1.288744037613344e+17, 1.288744037652408e+17, 1.288744037693032e+17, 1.288744037732095e+17, 1.288744037772719e+17, 1.288744037813345e+17, 1.288744037852408e+17, 1.288744037893032e+17, 1.288744037932096e+17, 1.288744037972719e+17, 1.288744038013345e+17, 1.288744038052407e+17, 1.288744038093032e+17, 1.288744038132095e+17, 1.288744038172719e+17, 1.288744038213345e+17, 1.288744038252407e+17, 1.288744038293033e+17, 1.288744038332095e+17, 1.288744038372719e+17, 1.288744038413345e+17, 1.288744038452407e+17, 1.288744038493032e+17, 1.288744038532095e+17, 1.288744038572719e+17, 1.288744038613345e+17, 1.288744038652407e+17, 1.288744038693033e+17, 1.288744038732095e+17, 1.288744038772721e+17, 1.288744038813345e+17, 1.288744038852407e+17, 1.288744038893033e+17, 1.288744038932095e+17, 1.288744038972719e+17, 1.288744039013345e+17, 1.288744039052407e+17, 1.288744039093033e+17, 1.288744039132095e+17, 1.288744039172721e+17, 1.288744039213345e+17, 1.288744039252407e+17, 1.288744039293033e+17, 1.288744039332095e+17, 1.288744039372721e+17, 1.288744039413345e+17, 1.288744039452407e+17, 1.288744039493033e+17, 1.288744039532095e+17, 1.288744039572721e+17, 1.288744039613344e+17, 1.288744039652408e+17, 1.288744039693033e+17, 1.288744039732095e+17, 1.288744039772721e+17, 1.288744039813344e+17, 1.288744039852407e+17, 1.288744039893032e+17, 1.288744039932095e+17, 1.288744039972721e+17, 1.288744040013345e+17, 1.288744040052408e+17, 1.288744040093032e+17, 1.288744040132095e+17, 1.288744040172719e+17, 1.288744040213344e+17, 1.288744040252408e+17, 1.288744040293032e+17, 1.288744040332095e+17, 1.288744040372719e+17, 1.288744040413345e+17, 1.288744040452407e+17, 1.288744040493033e+17, 1.288744040532096e+17, 1.288744040572719e+17, 1.288744040613345e+17, 1.288744040652407e+17, 1.288744040693032e+17, 1.288744040732095e+17, 1.288744040772719e+17, 1.288744040813345e+17, 1.288744040852407e+17, 1.288744040893033e+17, 1.288744040932095e+17, 1.288744040972719e+17, 1.288744041013345e+17, 1.288744041052407e+17, 1.288744041093032e+17, 1.288744041132095e+17, 1.288744041172719e+17, 1.288744041213345e+17, 1.288744041252407e+17, 1.288744041293033e+17, 1.288744041332095e+17, 1.288744041372721e+17, 1.288744041413345e+17, 1.288744041452407e+17, 1.288744041493033e+17, 1.288744041532095e+17, 1.288744041572719e+17, 1.288744041613345e+17, 1.288744041652407e+17, 1.288744041693033e+17, 1.288744041732095e+17, 1.288744041772721e+17, 1.288744041813345e+17, 1.288744041852407e+17, 1.288744041893033e+17, 1.288744041932095e+17, 1.288744041972721e+17, 1.288744042013345e+17, 1.288744042052407e+17, 1.288744042093033e+17, 1.288744042132095e+17, 1.288744042172721e+17, 1.288744042213344e+17, 1.288744042252408e+17, 1.288744042293033e+17, 1.288744042332095e+17, 1.288744042372721e+17, 1.288744042413344e+17, 1.288744042452407e+17, 1.288744042493032e+17, 1.288744042532095e+17, 1.288744042572721e+17, 1.288744042613345e+17, 1.288744042652408e+17, 1.288744042693032e+17, 1.288744042732096e+17, 1.288744042772719e+17, 1.288744042813344e+17, 1.288744042852408e+17, 1.288744042893032e+17, 1.288744042932095e+17, 1.288744042972719e+17, 1.288744043013345e+17, 1.288744043052407e+17, 1.288744043093033e+17, 1.288744043132096e+17, 1.288744043172719e+17, 1.288744043213345e+17, 1.288744043252407e+17, 1.288744043293032e+17, 1.288744043332095e+17, 1.288744043372719e+17, 1.288744043413345e+17, 1.288744043452407e+17, 1.288744043493033e+17, 1.288744043532095e+17, 1.288744043572719e+17, 1.288744043613345e+17, 1.288744043652407e+17, 1.288744043693033e+17, 1.288744043732095e+17, 1.288744043772719e+17, 1.288744043813345e+17, 1.288744043852407e+17, 1.288744043893033e+17, 1.288744043932095e+17, 1.288744043972721e+17, 1.288744044013345e+17, 1.288744044052407e+17, 1.288744044093033e+17, 1.288744044132095e+17, 1.288744044172719e+17, 1.288744044213345e+17, 1.288744044252407e+17, 1.288744044293033e+17, 1.288744044332095e+17, 1.288744044372721e+17, 1.288744044413345e+17, 1.288744044452407e+17, 1.288744044493033e+17, 1.288744044532095e+17, 1.288744044572721e+17, 1.288744044613345e+17, 1.288744044652407e+17, 1.288744044693033e+17, 1.288744044732095e+17, 1.288744044772721e+17, 1.288744044813344e+17, 1.288744044852408e+17, 1.288744044893033e+17, 1.288744044932095e+17, 1.288744044972721e+17, 1.288744045013344e+17, 1.288744045052407e+17, 1.288744045093032e+17, 1.288744045132095e+17, 1.288744045172721e+17, 1.288744045213345e+17, 1.288744045252408e+17, 1.288744045293032e+17, 1.288744045332096e+17, 1.288744045372719e+17, 1.288744045413344e+17, 1.288744045452408e+17, 1.288744045493032e+17, 1.288744045532095e+17, 1.288744045572719e+17, 1.288744045613345e+17, 1.288744045652407e+17, 1.288744045693033e+17, 1.288744045732096e+17, 1.288744045772719e+17, 1.288744045813345e+17, 1.288744045852407e+17, 1.288744045893032e+17, 1.288744045932095e+17, 1.288744045972719e+17, 1.288744046013345e+17, 1.288744046052407e+17, 1.288744046093033e+17, 1.288744046132095e+17, 1.288744046172719e+17, 1.288744046213345e+17, 1.288744046252407e+17, 1.288744046293033e+17, 1.288744046332095e+17, 1.288744046372719e+17, 1.288744046413345e+17, 1.288744046452407e+17, 1.288744046493033e+17, 1.288744046532095e+17, 1.288744046572721e+17, 1.288744046613345e+17, 1.288744046652407e+17, 1.288744046693033e+17, 1.288744046732095e+17, 1.288744046772719e+17, 1.288744046813345e+17, 1.288744046852407e+17, 1.288744046893033e+17, 1.288744046932095e+17, 1.288744046972721e+17, 1.288744047013345e+17, 1.288744047052407e+17, 1.288744047093033e+17, 1.288744047132095e+17, 1.288744047172721e+17, 1.288744047213345e+17, 1.288744047252407e+17, 1.288744047293033e+17, 1.288744047332095e+17, 1.288744047372721e+17, 1.288744047413345e+17, 1.288744047452408e+17, 1.288744047493033e+17, 1.288744047532095e+17, 1.288744047572721e+17, 1.288744047613344e+17, 1.288744047652407e+17, 1.288744047693032e+17, 1.288744047732095e+17, 1.288744047772721e+17, 1.288744047813345e+17, 1.288744047852408e+17, 1.288744047893032e+17, 1.288744047932096e+17, 1.288744047972719e+17, 1.288744048013344e+17, 1.288744048052408e+17, 1.288744048093032e+17, 1.288744048132095e+17, 1.288744048172719e+17, 1.288744048213345e+17, 1.288744048252407e+17, 1.288744048293033e+17, 1.288744048332096e+17, 1.288744048372719e+17, 1.288744048413345e+17, 1.288744048452407e+17, 1.288744048493032e+17, 1.288744048532095e+17, 1.288744048572719e+17, 1.288744048613345e+17, 1.288744048652407e+17, 1.288744048693033e+17, 1.288744048732095e+17, 1.288744048772719e+17, 1.288744048813345e+17, 1.288744048852407e+17, 1.288744048893033e+17, 1.288744048932095e+17, 1.288744048972719e+17, 1.288744049013345e+17, 1.288744049052407e+17, 1.288744049093033e+17, 1.288744049132095e+17, 1.288744049172721e+17, 1.288744049213345e+17, 1.288744049252407e+17, 1.288744049293033e+17, 1.288744049332095e+17, 1.288744049372719e+17, 1.288744049413345e+17, 1.288744049452407e+17, 1.288744049493033e+17, 1.288744049532095e+17, 1.288744049572721e+17, 1.288744049613345e+17, 1.288744049652408e+17, 1.288744049693033e+17, 1.288744049732095e+17, 1.288744049772721e+17, 1.288744049813344e+17, 1.288744049852407e+17, 1.288744049893033e+17, 1.288744049932095e+17, 1.288744049972721e+17, 1.288744050013345e+17, 1.288744050052408e+17, 1.288744050093032e+17, 1.288744050132095e+17, 1.288744050172721e+17, 1.288744050213344e+17, 1.288744050252408e+17, 1.288744050293032e+17, 1.288744050332095e+17, 1.288744050372719e+17, 1.288744050413345e+17, 1.288744050452408e+17, 1.288744050493032e+17, 1.288744050532096e+17, 1.288744050572719e+17, 1.288744050613345e+17, 1.288744050652407e+17, 1.288744050693032e+17, 1.288744050732095e+17, 1.288744050772719e+17, 1.288744050813345e+17, 1.288744050852407e+17, 1.288744050893033e+17, 1.288744050932095e+17, 1.288744050972719e+17, 1.288744051013345e+17, 1.288744051052407e+17, 1.288744051093032e+17, 1.288744051132095e+17, 1.288744051172719e+17, 1.288744051213345e+17, 1.288744051252407e+17, 1.288744051293033e+17, 1.288744051332095e+17, 1.288744051372719e+17, 1.288744051413345e+17, 1.288744051452407e+17, 1.288744051493033e+17, 1.288744051532095e+17, 1.288744051572719e+17, 1.288744051613345e+17, 1.288744051652407e+17, 1.288744051693033e+17, 1.288744051732095e+17, 1.288744051772721e+17, 1.288744051813345e+17, 1.288744051852407e+17, 1.288744051893033e+17, 1.288744051932095e+17, 1.288744051972719e+17, 1.288744052013345e+17, 1.288744052052407e+17, 1.288744052093033e+17, 1.288744052132095e+17, 1.288744052172721e+17, 1.288744052213345e+17, 1.288744052252408e+17, 1.288744052293033e+17, 1.288744052332095e+17, 1.288744052372721e+17, 1.288744052413344e+17, 1.288744052452407e+17, 1.288744052493033e+17, 1.288744052532095e+17, 1.288744052572721e+17, 1.288744052613345e+17, 1.288744052652408e+17, 1.288744052693032e+17, 1.288744052732095e+17, 1.288744052772721e+17, 1.288744052813344e+17, 1.288744052852408e+17, 1.288744052893032e+17, 1.288744052932095e+17, 1.288744052972719e+17, 1.288744053013345e+17, 1.288744053052408e+17, 1.288744053093032e+17, 1.288744053132096e+17, 1.288744053172719e+17, 1.288744053213345e+17, 1.288744053252407e+17, 1.288744053293032e+17, 1.288744053332095e+17, 1.288744053372719e+17, 1.288744053413345e+17, 1.288744053452407e+17, 1.288744053493033e+17, 1.288744053532095e+17, 1.288744053572719e+17, 1.288744053613345e+17, 1.288744053652407e+17, 1.288744053693032e+17, 1.288744053732095e+17, 1.288744053772719e+17, 1.288744053813345e+17, 1.288744053852407e+17, 1.288744053893033e+17, 1.288744053932095e+17, 1.288744053972721e+17, 1.288744054013345e+17, 1.288744054052407e+17, 1.288744054093033e+17, 1.288744054132095e+17, 1.288744054172719e+17, 1.288744054213345e+17, 1.288744054252407e+17, 1.288744054293033e+17, 1.288744054332095e+17, 1.288744054372721e+17, 1.288744054413345e+17, 1.288744054452407e+17, 1.288744054493033e+17, 1.288744054532095e+17, 1.288744054572719e+17, 1.288744054613345e+17, 1.288744054652407e+17, 1.288744054693033e+17, 1.288744054732095e+17, 1.288744054772721e+17, 1.288744054813345e+17, 1.288744054852408e+17, 1.288744054893033e+17, 1.288744054932095e+17, 1.288744054972721e+17, 1.288744055013344e+17, 1.288744055052407e+17, 1.288744055093033e+17, 1.288744055132095e+17, 1.288744055172721e+17, 1.288744055213345e+17, 1.288744055252408e+17, 1.288744055293032e+17, 1.288744055332095e+17, 1.288744055372721e+17, 1.288744055413344e+17, 1.288744055452408e+17, 1.288744055493032e+17, 1.288744055532095e+17, 1.288744055572719e+17, 1.288744055613345e+17, 1.288744055652408e+17, 1.288744055693032e+17, 1.288744055732096e+17, 1.288744055772719e+17, 1.288744055813345e+17, 1.288744055852407e+17, 1.288744055893032e+17, 1.288744055932095e+17, 1.288744055972719e+17, 1.288744056013345e+17, 1.288744056052407e+17, 1.288744056093033e+17, 1.288744056132095e+17, 1.288744056172719e+17, 1.288744056213345e+17, 1.288744056252407e+17, 1.288744056293032e+17, 1.288744056332095e+17, 1.288744056372719e+17, 1.288744056413345e+17, 1.288744056452407e+17, 1.288744056493033e+17, 1.288744056532095e+17, 1.288744056572721e+17, 1.288744056613345e+17, 1.288744056652407e+17, 1.288744056693033e+17, 1.288744056732095e+17, 1.288744056772719e+17, 1.288744056813345e+17, 1.288744056852407e+17, 1.288744056893033e+17, 1.288744056932095e+17, 1.288744056972721e+17, 1.288744057013345e+17, 1.288744057052407e+17, 1.288744057093033e+17, 1.288744057132095e+17, 1.288744057172721e+17, 1.288744057213345e+17, 1.288744057252407e+17, 1.288744057293033e+17, 1.288744057332095e+17, 1.288744057372721e+17, 1.288744057413345e+17, 1.288744057452408e+17, 1.288744057493033e+17, 1.288744057532095e+17, 1.288744057572721e+17, 1.288744057613344e+17, 1.288744057652407e+17, 1.288744057693033e+17, 1.288744057732095e+17, 1.288744057772721e+17, 1.288744057813345e+17, 1.288744057852408e+17, 1.288744057893032e+17, 1.288744057932095e+17, 1.288744057972721e+17, 1.288744058013344e+17, 1.288744058052408e+17, 1.288744058093032e+17, 1.288744058132095e+17, 1.288744058172719e+17, 1.288744058213345e+17, 1.288744058252408e+17, 1.288744058293032e+17, 1.288744058332096e+17, 1.288744058372719e+17, 1.288744058413345e+17, 1.288744058452407e+17, 1.288744058493032e+17, 1.288744058532095e+17, 1.288744058572719e+17, 1.288744058613345e+17, 1.288744058652407e+17, 1.288744058693033e+17, 1.288744058732095e+17, 1.288744058772719e+17, 1.288744058813345e+17, 1.288744058852407e+17, 1.288744058893032e+17, 1.288744058932095e+17, 1.288744058972719e+17, 1.288744059013345e+17, 1.288744059052407e+17, 1.288744059093033e+17, 1.288744059132095e+17, 1.288744059172721e+17, 1.288744059213345e+17, 1.288744059252407e+17, 1.288744059293033e+17, 1.288744059332095e+17, 1.288744059372719e+17, 1.288744059413345e+17, 1.288744059452407e+17, 1.288744059493033e+17, 1.288744059532095e+17, 1.288744059572721e+17, 1.288744059613345e+17, 1.288744059652407e+17, 1.288744059693033e+17, 1.288744059732095e+17, 1.288744059772721e+17, 1.288744059813345e+17, 1.288744059852407e+17, 1.288744059893033e+17, 1.288744059932095e+17, 1.288744059972721e+17, 1.288744060013344e+17, 1.288744060052408e+17, 1.288744060093033e+17, 1.288744060132095e+17, 1.288744060172721e+17, 1.288744060213344e+17, 1.288744060252407e+17, 1.288744060293032e+17, 1.288744060332095e+17, 1.288744060372721e+17, 1.288744060413345e+17, 1.288744060452408e+17, 1.288744060493032e+17, 1.288744060532096e+17, 1.288744060572719e+17, 1.288744060613344e+17, 1.288744060652408e+17, 1.288744060693032e+17, 1.288744060732095e+17, 1.288744060772719e+17, 1.288744060813345e+17, 1.288744060852407e+17, 1.288744060893033e+17, 1.288744060932096e+17, 1.288744060972719e+17, 1.288744061013345e+17, 1.288744061052407e+17, 1.288744061093032e+17, 1.288744061132095e+17, 1.288744061172719e+17, 1.288744061213345e+17, 1.288744061252407e+17, 1.288744061293033e+17, 1.288744061332095e+17, 1.288744061372719e+17, 1.288744061413345e+17, 1.288744061452407e+17, 1.288744061493032e+17, 1.288744061532095e+17, 1.288744061572719e+17, 1.288744061613345e+17, 1.288744061652407e+17, 1.288744061693033e+17, 1.288744061732095e+17, 1.288744061772721e+17, 1.288744061813345e+17, 1.288744061852407e+17, 1.288744061893033e+17, 1.288744061932095e+17, 1.288744061972719e+17, 1.288744062013345e+17, 1.288744062052407e+17, 1.288744062093033e+17, 1.288744062132095e+17, 1.288744062172721e+17, 1.288744062213345e+17, 1.288744062252407e+17, 1.288744062293033e+17, 1.288744062332095e+17, 1.288744062372721e+17, 1.288744062413345e+17, 1.288744062452407e+17, 1.288744062493033e+17, 1.288744062532095e+17, 1.288744062572721e+17, 1.288744062613344e+17, 1.288744062652408e+17, 1.288744062693033e+17, 1.288744062732095e+17, 1.288744062772721e+17, 1.288744062813344e+17, 1.288744062852407e+17, 1.288744062893032e+17, 1.288744062932095e+17, 1.288744062972721e+17, 1.288744063013345e+17, 1.288744063052408e+17, 1.288744063093032e+17, 1.288744063132096e+17, 1.288744063172719e+17, 1.288744063213344e+17, 1.288744063252408e+17, 1.288744063293032e+17, 1.288744063332095e+17, 1.288744063372719e+17, 1.288744063413345e+17, 1.288744063452407e+17, 1.288744063493033e+17, 1.288744063532096e+17, 1.288744063572719e+17, 1.288744063613345e+17, 1.288744063652407e+17, 1.288744063693032e+17, 1.288744063732095e+17, 1.288744063772719e+17, 1.288744063813345e+17, 1.288744063852407e+17, 1.288744063893033e+17, 1.288744063932095e+17, 1.288744063972719e+17, 1.288744064013345e+17, 1.288744064052407e+17, 1.288744064093033e+17, 1.288744064132095e+17, 1.288744064172719e+17, 1.288744064213345e+17, 1.288744064252407e+17, 1.288744064293033e+17, 1.288744064332095e+17, 1.288744064372721e+17, 1.288744064413345e+17, 1.288744064452407e+17, 1.288744064493033e+17, 1.288744064532095e+17, 1.288744064572719e+17, 1.288744064613345e+17, 1.288744064652407e+17, 1.288744064693033e+17, 1.288744064732095e+17, 1.288744064772721e+17, 1.288744064813345e+17, 1.288744064852407e+17, 1.288744064893033e+17, 1.288744064932095e+17, 1.288744064972721e+17, 1.288744065013345e+17, 1.288744065052407e+17, 1.288744065093033e+17, 1.288744065132095e+17, 1.288744065172721e+17, 1.288744065213344e+17, 1.288744065252408e+17, 1.288744065293033e+17, 1.288744065332095e+17, 1.288744065372721e+17, 1.288744065413344e+17, 1.288744065452407e+17, 1.288744065493032e+17, 1.288744065532095e+17, 1.288744065572721e+17, 1.288744065613345e+17, 1.288744065652408e+17, 1.288744065693032e+17, 1.288744065732096e+17, 1.288744065772719e+17, 1.288744065813344e+17, 1.288744065852408e+17, 1.288744065893032e+17, 1.288744065932095e+17, 1.288744065972719e+17, 1.288744066013345e+17, 1.288744066052407e+17, 1.288744066093033e+17, 1.288744066132096e+17, 1.288744066172719e+17, 1.288744066213345e+17, 1.288744066252407e+17, 1.288744066293032e+17, 1.288744066332095e+17, 1.288744066372719e+17, 1.288744066413345e+17, 1.288744066452407e+17, 1.288744066493033e+17, 1.288744066532095e+17, 1.288744066572719e+17, 1.288744066613345e+17, 1.288744066652407e+17, 1.288744066693033e+17, 1.288744066732095e+17, 1.288744066772719e+17, 1.288744066813345e+17, 1.288744066852407e+17, 1.288744066893033e+17, 1.288744066932095e+17, 1.288744066972721e+17, 1.288744067013345e+17, 1.288744067052407e+17, 1.288744067093033e+17, 1.288744067132095e+17, 1.288744067172719e+17, 1.288744067213345e+17, 1.288744067252407e+17, 1.288744067293033e+17, 1.288744067332095e+17, 1.288744067372721e+17, 1.288744067413345e+17, 1.288744067452408e+17, 1.288744067493033e+17, 1.288744067532095e+17, 1.288744067572721e+17, 1.288744067613344e+17, 1.288744067652407e+17, 1.288744067693033e+17, 1.288744067732095e+17, 1.288744067772721e+17, 1.288744067813345e+17, 1.288744067852408e+17, 1.288744067893032e+17, 1.288744067932095e+17, 1.288744067972721e+17, 1.288744068013344e+17, 1.288744068052407e+17, 1.288744068093032e+17, 1.288744068132095e+17, 1.288744068172721e+17, 1.288744068213345e+17, 1.288744068252408e+17, 1.288744068293032e+17, 1.288744068332096e+17, 1.288744068372719e+17, 1.288744068413345e+17, 1.288744068452408e+17, 1.288744068493032e+17, 1.288744068532095e+17, 1.288744068572719e+17, 1.288744068613345e+17, 1.288744068652407e+17, 1.288744068693033e+17, 1.288744068732096e+17, 1.288744068772719e+17, 1.288744068813345e+17, 1.288744068852407e+17, 1.288744068893032e+17, 1.288744068932095e+17, 1.288744068972719e+17, 1.288744069013345e+17, 1.288744069052407e+17, 1.288744069093033e+17, 1.288744069132095e+17, 1.288744069172719e+17, 1.288744069213345e+17, 1.288744069252407e+17, 1.288744069293033e+17, 1.288744069332095e+17, 1.288744069372719e+17, 1.288744069413345e+17, 1.288744069452407e+17, 1.288744069493033e+17, 1.288744069532095e+17, 1.288744069572721e+17, 1.288744069613345e+17, 1.288744069652407e+17, 1.288744069693033e+17, 1.288744069732095e+17, 1.288744069772719e+17, 1.288744069813345e+17, 1.288744069852407e+17, 1.288744069893033e+17, 1.288744069932095e+17, 1.288744069972721e+17, 1.288744070013345e+17, 1.288744070052408e+17, 1.288744070093033e+17, 1.288744070132095e+17, 1.288744070172721e+17, 1.288744070213344e+17, 1.288744070252407e+17, 1.288744070293033e+17, 1.288744070332095e+17, 1.288744070372721e+17, 1.288744070413345e+17, 1.288744070452408e+17, 1.288744070493032e+17, 1.288744070532095e+17, 1.288744070572721e+17, 1.288744070613344e+17, 1.288744070652408e+17, 1.288744070693032e+17, 1.288744070732095e+17, 1.288744070772719e+17, 1.288744070813345e+17, 1.288744070852408e+17, 1.288744070893032e+17, 1.288744070932096e+17, 1.288744070972719e+17, 1.288744071013345e+17, 1.288744071052407e+17, 1.288744071093032e+17, 1.288744071132095e+17, 1.288744071172719e+17, 1.288744071213345e+17, 1.288744071252407e+17, 1.288744071293033e+17, 1.288744071332095e+17, 1.288744071372719e+17, 1.288744071413345e+17, 1.288744071452407e+17, 1.288744071493032e+17, 1.288744071532095e+17, 1.288744071572719e+17, 1.288744071613345e+17, 1.288744071652407e+17, 1.288744071693033e+17, 1.288744071732095e+17, 1.288744071772719e+17, 1.288744071813345e+17, 1.288744071852407e+17, 1.288744071893033e+17, 1.288744071932095e+17, 1.288744071972719e+17, 1.288744072013345e+17, 1.288744072052407e+17, 1.288744072093033e+17, 1.288744072132095e+17, 1.288744072172721e+17, 1.288744072213345e+17, 1.288744072252407e+17, 1.288744072293033e+17, 1.288744072332095e+17, 1.288744072372719e+17, 1.288744072413345e+17, 1.288744072452407e+17, 1.288744072493033e+17, 1.288744072532095e+17, 1.288744072572721e+17, 1.288744072613345e+17, 1.288744072652408e+17, 1.288744072693033e+17, 1.288744072732095e+17, 1.288744072772721e+17, 1.288744072813344e+17, 1.288744072852407e+17, 1.288744072893033e+17, 1.288744072932095e+17, 1.288744072972721e+17, 1.288744073013345e+17, 1.288744073052408e+17, 1.288744073093032e+17, 1.288744073132095e+17, 1.288744073172721e+17, 1.288744073213344e+17, 1.288744073252408e+17, 1.288744073293032e+17, 1.288744073332095e+17, 1.288744073372719e+17, 1.288744073413345e+17, 1.288744073452408e+17, 1.288744073493032e+17, 1.288744073532096e+17, 1.288744073572719e+17, 1.288744073613345e+17, 1.288744073652407e+17, 1.288744073693032e+17, 1.288744073732095e+17, 1.288744073772719e+17, 1.288744073813345e+17, 1.288744073852407e+17, 1.288744073893033e+17, 1.288744073932095e+17, 1.288744073972719e+17, 1.288744074013345e+17, 1.288744074052407e+17, 1.288744074093032e+17, 1.288744074132095e+17, 1.288744074172719e+17, 1.288744074213345e+17, 1.288744074252407e+17, 1.288744074293033e+17, 1.288744074332095e+17, 1.288744074372721e+17, 1.288744074413345e+17, 1.288744074452407e+17, 1.288744074493033e+17, 1.288744074532095e+17, 1.288744074572719e+17, 1.288744074613345e+17, 1.288744074652407e+17, 1.288744074693033e+17, 1.288744074732095e+17, 1.288744074772721e+17, 1.288744074813345e+17, 1.288744074852407e+17, 1.288744074893033e+17, 1.288744074932095e+17, 1.288744074972721e+17, 1.288744075013345e+17, 1.288744075052407e+17, 1.288744075093033e+17, 1.288744075132095e+17, 1.288744075172721e+17, 1.288744075213345e+17, 1.288744075252408e+17, 1.288744075293033e+17, 1.288744075332095e+17, 1.288744075372721e+17, 1.288744075413344e+17, 1.288744075452407e+17, 1.288744075493033e+17, 1.288744075532095e+17, 1.288744075572721e+17, 1.288744075613345e+17, 1.288744075652408e+17, 1.288744075693032e+17, 1.288744075732095e+17, 1.288744075772721e+17, 1.288744075813344e+17, 1.288744075852408e+17, 1.288744075893032e+17, 1.288744075932095e+17, 1.288744075972719e+17, 1.288744076013345e+17, 1.288744076052408e+17, 1.288744076093032e+17, 1.288744076132096e+17, 1.288744076172719e+17, 1.288744076213345e+17, 1.288744076252407e+17, 1.288744076293032e+17, 1.288744076332095e+17, 1.288744076372719e+17, 1.288744076413345e+17, 1.288744076452407e+17, 1.288744076493033e+17, 1.288744076532095e+17, 1.288744076572719e+17, 1.288744076613345e+17, 1.288744076652407e+17, 1.288744076693032e+17, 1.288744076732095e+17, 1.288744076772719e+17, 1.288744076813345e+17, 1.288744076852407e+17, 1.288744076893033e+17, 1.288744076932095e+17, 1.288744076972721e+17, 1.288744077013345e+17, 1.288744077052407e+17, 1.288744077093033e+17, 1.288744077132095e+17, 1.288744077172719e+17, 1.288744077213345e+17, 1.288744077252407e+17, 1.288744077293033e+17, 1.288744077332095e+17, 1.288744077372721e+17, 1.288744077413345e+17, 1.288744077452407e+17, 1.288744077493033e+17, 1.288744077532095e+17, 1.288744077572721e+17, 1.288744077613345e+17, 1.288744077652407e+17, 1.288744077693033e+17, 1.288744077732095e+17, 1.288744077772721e+17, 1.288744077813344e+17, 1.288744077852408e+17, 1.288744077893033e+17, 1.288744077932095e+17, 1.288744077972721e+17, 1.288744078013344e+17, 1.288744078052407e+17, 1.288744078093032e+17, 1.288744078132095e+17, 1.288744078172721e+17, 1.288744078213345e+17, 1.288744078252408e+17, 1.288744078293032e+17, 1.288744078332095e+17, 1.288744078372719e+17, 1.288744078413344e+17, 1.288744078452408e+17, 1.288744078493032e+17, 1.288744078532095e+17, 1.288744078572719e+17, 1.288744078613345e+17, 1.288744078652407e+17, 1.288744078693032e+17, 1.288744078732096e+17, 1.288744078772719e+17, 1.288744078813345e+17, 1.288744078852407e+17, 1.288744078893032e+17, 1.288744078932095e+17, 1.288744078972719e+17, 1.288744079013345e+17, 1.288744079052407e+17, 1.288744079093033e+17, 1.288744079132095e+17, 1.288744079172719e+17, 1.288744079213345e+17, 1.288744079252407e+17, 1.288744079293032e+17, 1.288744079332095e+17, 1.288744079372719e+17, 1.288744079413345e+17, 1.288744079452407e+17, 1.288744079493033e+17, 1.288744079532095e+17, 1.288744079572721e+17, 1.288744079613345e+17, 1.288744079652407e+17, 1.288744079693033e+17, 1.288744079732095e+17, 1.288744079772719e+17, 1.288744079813345e+17, 1.288744079852407e+17, 1.288744079893033e+17, 1.288744079932095e+17, 1.288744079972721e+17, 1.288744080013345e+17, 1.288744080052407e+17, 1.288744080093033e+17, 1.288744080132095e+17, 1.288744080172721e+17, 1.288744080213345e+17, 1.288744080252407e+17, 1.288744080293033e+17, 1.288744080332095e+17, 1.288744080372721e+17, 1.288744080413344e+17, 1.288744080452408e+17, 1.288744080493033e+17, 1.288744080532095e+17, 1.288744080572721e+17, 1.288744080613344e+17, 1.288744080652407e+17, 1.288744080693032e+17, 1.288744080732095e+17, 1.288744080772721e+17, 1.288744080813345e+17, 1.288744080852408e+17, 1.288744080893032e+17, 1.288744080932096e+17, 1.288744080972719e+17, 1.288744081013344e+17, 1.288744081052408e+17, 1.288744081093032e+17, 1.288744081132095e+17, 1.288744081172719e+17, 1.288744081213345e+17, 1.288744081252407e+17, 1.288744081293033e+17, 1.288744081332096e+17, 1.288744081372719e+17, 1.288744081413345e+17, 1.288744081452407e+17, 1.288744081493032e+17, 1.288744081532095e+17, 1.288744081572719e+17, 1.288744081613345e+17, 1.288744081652407e+17, 1.288744081693033e+17, 1.288744081732095e+17, 1.288744081772719e+17, 1.288744081813345e+17, 1.288744081852407e+17, 1.288744081893033e+17, 1.288744081932095e+17, 1.288744081972719e+17, 1.288744082013345e+17, 1.288744082052407e+17, 1.288744082093033e+17, 1.288744082132095e+17, 1.288744082172721e+17, 1.288744082213345e+17, 1.288744082252407e+17, 1.288744082293033e+17, 1.288744082332095e+17, 1.288744082372719e+17, 1.288744082413345e+17, 1.288744082452407e+17, 1.288744082493033e+17, 1.288744082532095e+17, 1.288744082572721e+17, 1.288744082613345e+17, 1.288744082652407e+17, 1.288744082693033e+17, 1.288744082732095e+17, 1.288744082772721e+17, 1.288744082813345e+17, 1.288744082852407e+17, 1.288744082893033e+17, 1.288744082932095e+17, 1.288744082972721e+17, 1.288744083013344e+17, 1.288744083052408e+17, 1.288744083093033e+17, 1.288744083132095e+17, 1.288744083172721e+17, 1.288744083213344e+17, 1.288744083252407e+17, 1.288744083293032e+17, 1.288744083332095e+17, 1.288744083372721e+17, 1.288744083413345e+17, 1.288744083452408e+17, 1.288744083493032e+17, 1.288744083532096e+17, 1.288744083572719e+17, 1.288744083613344e+17, 1.288744083652408e+17, 1.288744083693032e+17, 1.288744083732095e+17, 1.288744083772719e+17, 1.288744083813345e+17, 1.288744083852407e+17, 1.288744083893033e+17, 1.288744083932096e+17, 1.288744083972719e+17, 1.288744084013345e+17, 1.288744084052407e+17, 1.288744084093032e+17, 1.288744084132095e+17, 1.288744084172719e+17, 1.288744084213345e+17, 1.288744084252407e+17, 1.288744084293033e+17, 1.288744084332095e+17, 1.288744084372719e+17, 1.288744084413345e+17, 1.288744084452407e+17, 1.288744084493033e+17, 1.288744084532095e+17, 1.288744084572719e+17, 1.288744084613345e+17, 1.288744084652407e+17, 1.288744084693033e+17, 1.288744084732095e+17, 1.288744084772721e+17, 1.288744084813345e+17, 1.288744084852407e+17, 1.288744084893033e+17, 1.288744084932095e+17, 1.288744084972719e+17, 1.288744085013345e+17, 1.288744085052407e+17, 1.288744085093033e+17, 1.288744085132095e+17, 1.288744085172721e+17, 1.288744085213345e+17, 1.288744085252407e+17, 1.288744085293033e+17, 1.288744085332095e+17, 1.288744085372721e+17, 1.288744085413345e+17, 1.288744085452407e+17, 1.288744085493033e+17, 1.288744085532095e+17, 1.288744085572721e+17, 1.288744085613345e+17, 1.288744085652408e+17, 1.288744085693033e+17, 1.288744085732095e+17, 1.288744085772721e+17, 1.288744085813344e+17, 1.288744085852407e+17, 1.288744085893032e+17, 1.288744085932095e+17, 1.288744085972721e+17, 1.288744086013345e+17, 1.288744086052408e+17, 1.288744086093032e+17, 1.288744086132096e+17, 1.288744086172719e+17, 1.288744086213344e+17, 1.288744086252408e+17, 1.288744086293032e+17, 1.288744086332095e+17, 1.288744086372719e+17, 1.288744086413345e+17, 1.288744086452407e+17, 1.288744086493033e+17, 1.288744086532096e+17, 1.288744086572719e+17, 1.288744086613345e+17, 1.288744086652407e+17, 1.288744086693032e+17, 1.288744086732095e+17, 1.288744086772719e+17, 1.288744086813345e+17, 1.288744086852407e+17, 1.288744086893033e+17, 1.288744086932095e+17, 1.288744086972719e+17, 1.288744087013345e+17, 1.288744087052407e+17, 1.288744087093033e+17, 1.288744087132095e+17, 1.288744087172719e+17, 1.288744087213345e+17, 1.288744087252407e+17, 1.288744087293033e+17, 1.288744087332095e+17, 1.288744087372721e+17, 1.288744087413345e+17, 1.288744087452407e+17, 1.288744087493033e+17, 1.288744087532095e+17, 1.288744087572719e+17, 1.288744087613345e+17, 1.288744087652407e+17, 1.288744087693033e+17, 1.288744087732095e+17, 1.288744087772721e+17, 1.288744087813345e+17, 1.288744087852408e+17, 1.288744087893033e+17, 1.288744087932095e+17, 1.288744087972721e+17, 1.288744088013344e+17, 1.288744088052407e+17, 1.288744088093033e+17, 1.288744088132095e+17, 1.288744088172721e+17, 1.288744088213345e+17, 1.288744088252408e+17, 1.288744088293032e+17, 1.288744088332095e+17, 1.288744088372721e+17, 1.288744088413344e+17, 1.288744088452408e+17, 1.288744088493032e+17, 1.288744088532095e+17, 1.288744088572719e+17, 1.288744088613345e+17, 1.288744088652408e+17, 1.288744088693032e+17, 1.288744088732096e+17, 1.288744088772719e+17, 1.288744088813345e+17, 1.288744088852407e+17, 1.288744088893032e+17, 1.288744088932095e+17, 1.288744088972719e+17, 1.288744089013345e+17, 1.288744089052407e+17, 1.288744089093033e+17, 1.288744089132095e+17, 1.288744089172719e+17, 1.288744089213345e+17, 1.288744089252407e+17, 1.288744089293032e+17, 1.288744089332095e+17, 1.288744089372719e+17, 1.288744089413345e+17, 1.288744089452407e+17, 1.288744089493033e+17, 1.288744089532095e+17, 1.288744089572719e+17, 1.288744089613345e+17, 1.288744089652407e+17, 1.288744089693033e+17, 1.288744089732095e+17, 1.288744089772719e+17, 1.288744089813345e+17, 1.288744089852407e+17, 1.288744089893033e+17, 1.288744089932095e+17, 1.288744089972721e+17, 1.288744090013345e+17, 1.288744090052407e+17, 1.288744090093033e+17, 1.288744090132095e+17, 1.288744090172719e+17, 1.288744090213345e+17, 1.288744090252407e+17, 1.288744090293033e+17, 1.288744090332095e+17, 1.288744090372721e+17, 1.288744090413345e+17, 1.288744090452408e+17, 1.288744090493033e+17, 1.288744090532095e+17, 1.288744090572721e+17, 1.288744090613344e+17, 1.288744090652407e+17, 1.288744090693033e+17, 1.288744090732095e+17, 1.288744090772721e+17, 1.288744090813345e+17, 1.288744090852408e+17, 1.288744090893032e+17, 1.288744090932095e+17, 1.288744090972721e+17, 1.288744091013344e+17, 1.288744091052408e+17, 1.288744091093032e+17, 1.288744091132095e+17, 1.288744091172719e+17, 1.288744091213345e+17, 1.288744091252408e+17, 1.288744091293032e+17, 1.288744091332096e+17, 1.288744091372719e+17, 1.288744091413345e+17, 1.288744091452407e+17, 1.288744091493032e+17, 1.288744091532095e+17, 1.288744091572719e+17, 1.288744091613345e+17, 1.288744091652407e+17, 1.288744091693033e+17, 1.288744091732095e+17, 1.288744091772719e+17, 1.288744091813345e+17, 1.288744091852407e+17, 1.288744091893032e+17, 1.288744091932095e+17, 1.288744091972719e+17, 1.288744092013345e+17, 1.288744092052407e+17, 1.288744092093033e+17, 1.288744092132095e+17, 1.288744092172721e+17, 1.288744092213345e+17, 1.288744092252407e+17, 1.288744092293033e+17, 1.288744092332095e+17, 1.288744092372719e+17, 1.288744092413345e+17, 1.288744092452407e+17, 1.288744092493033e+17, 1.288744092532095e+17, 1.288744092572721e+17, 1.288744092613345e+17, 1.288744092652407e+17, 1.288744092693033e+17, 1.288744092732095e+17, 1.288744092772719e+17, 1.288744092813345e+17, 1.288744092852407e+17, 1.288744092893033e+17, 1.288744092932095e+17, 1.288744092972721e+17, 1.288744093013345e+17, 1.288744093052408e+17, 1.288744093093033e+17, 1.288744093132095e+17, 1.288744093172721e+17, 1.288744093213344e+17, 1.288744093252407e+17, 1.288744093293033e+17, 1.288744093332095e+17, 1.288744093372721e+17, 1.288744093413345e+17, 1.288744093452408e+17, 1.288744093493032e+17, 1.288744093532095e+17, 1.288744093572721e+17, 1.288744093613344e+17, 1.288744093652408e+17, 1.288744093693032e+17, 1.288744093732095e+17, 1.288744093772719e+17, 1.288744093813345e+17, 1.288744093852408e+17, 1.288744093893032e+17, 1.288744093932096e+17, 1.288744093972719e+17, 1.288744094013345e+17, 1.288744094052407e+17, 1.288744094093032e+17, 1.288744094132095e+17, 1.288744094172719e+17, 1.288744094213345e+17, 1.288744094252407e+17, 1.288744094293033e+17, 1.288744094332095e+17, 1.288744094372719e+17, 1.288744094413345e+17, 1.288744094452407e+17, 1.288744094493032e+17, 1.288744094532095e+17, 1.288744094572719e+17, 1.288744094613345e+17, 1.288744094652407e+17, 1.288744094693033e+17, 1.288744094732095e+17, 1.288744094772721e+17, 1.288744094813345e+17, 1.288744094852407e+17, 1.288744094893033e+17, 1.288744094932095e+17, 1.288744094972719e+17, 1.288744095013345e+17, 1.288744095052407e+17, 1.288744095093033e+17, 1.288744095132095e+17, 1.288744095172721e+17, 1.288744095213345e+17, 1.288744095252407e+17, 1.288744095293033e+17, 1.288744095332095e+17, 1.288744095372721e+17, 1.288744095413345e+17, 1.288744095452407e+17, 1.288744095493033e+17, 1.288744095532095e+17, 1.288744095572721e+17, 1.288744095613345e+17, 1.288744095652408e+17, 1.288744095693033e+17, 1.288744095732095e+17, 1.288744095772721e+17, 1.288744095813344e+17, 1.288744095852407e+17, 1.288744095893033e+17, 1.288744095932095e+17, 1.288744095972721e+17, 1.288744096013345e+17, 1.288744096052408e+17, 1.288744096093032e+17, 1.288744096132095e+17, 1.288744096172721e+17, 1.288744096213344e+17, 1.288744096252408e+17, 1.288744096293032e+17, 1.288744096332095e+17, 1.288744096372719e+17, 1.288744096413345e+17, 1.288744096452408e+17, 1.288744096493032e+17, 1.288744096532096e+17, 1.288744096572719e+17, 1.288744096613345e+17, 1.288744096652407e+17, 1.288744096693032e+17, 1.288744096732095e+17, 1.288744096772719e+17, 1.288744096813345e+17, 1.288744096852407e+17, 1.288744096893033e+17, 1.288744096932095e+17, 1.288744096972719e+17, 1.288744097013345e+17, 1.288744097052407e+17, 1.288744097093032e+17, 1.288744097132095e+17, 1.288744097172719e+17, 1.288744097213345e+17, 1.288744097252407e+17, 1.288744097293033e+17, 1.288744097332095e+17, 1.288744097372721e+17, 1.288744097413345e+17, 1.288744097452407e+17, 1.288744097493033e+17, 1.288744097532095e+17, 1.288744097572719e+17, 1.288744097613345e+17, 1.288744097652407e+17, 1.288744097693033e+17, 1.288744097732095e+17, 1.288744097772721e+17, 1.288744097813345e+17, 1.288744097852407e+17, 1.288744097893033e+17, 1.288744097932095e+17, 1.288744097972721e+17, 1.288744098013345e+17, 1.288744098052407e+17, 1.288744098093033e+17, 1.288744098132095e+17, 1.288744098172721e+17, 1.288744098213344e+17, 1.288744098252408e+17, 1.288744098293033e+17, 1.288744098332095e+17, 1.288744098372721e+17, 1.288744098413344e+17, 1.288744098452407e+17, 1.288744098493032e+17, 1.288744098532095e+17, 1.288744098572721e+17, 1.288744098613345e+17, 1.288744098652408e+17, 1.288744098693032e+17, 1.288744098732095e+17, 1.288744098772719e+17, 1.288744098813344e+17, 1.288744098852408e+17, 1.288744098893032e+17, 1.288744098932095e+17, 1.288744098972719e+17, 1.288744099013345e+17, 1.288744099052407e+17, 1.288744099093033e+17, 1.288744099132096e+17, 1.288744099172719e+17, 1.288744099213345e+17, 1.288744099252407e+17, 1.288744099293032e+17, 1.288744099332095e+17, 1.288744099372719e+17, 1.288744099413345e+17, 1.288744099452407e+17, 1.288744099493033e+17, 1.288744099532095e+17, 1.288744099572719e+17, 1.288744099613345e+17, 1.288744099652407e+17, 1.288744099693032e+17, 1.288744099732095e+17, 1.288744099772719e+17, 1.288744099813345e+17, 1.288744099852407e+17, 1.288744099893033e+17, 1.288744099932095e+17, 1.288744099972721e+17, 1.288744100013345e+17, 1.288744100052407e+17, 1.288744100093033e+17, 1.288744100132095e+17, 1.288744100172719e+17, 1.288744100213345e+17, 1.288744100252407e+17, 1.288744100293033e+17, 1.288744100332095e+17, 1.288744100372721e+17, 1.288744100413345e+17, 1.288744100452407e+17, 1.288744100493033e+17, 1.288744100532095e+17, 1.288744100572721e+17, 1.288744100613345e+17, 1.288744100652407e+17, 1.288744100693033e+17, 1.288744100732095e+17, 1.288744100772721e+17, 1.288744100813344e+17, 1.288744100852408e+17, 1.288744100893033e+17, 1.288744100932095e+17, 1.288744100972721e+17, 1.288744101013344e+17, 1.288744101052407e+17, 1.288744101093032e+17, 1.288744101132095e+17, 1.288744101172721e+17, 1.288744101213345e+17, 1.288744101252408e+17, 1.288744101293032e+17, 1.288744101332096e+17, 1.288744101372719e+17, 1.288744101413344e+17, 1.288744101452408e+17, 1.288744101493032e+17, 1.288744101532095e+17, 1.288744101572719e+17, 1.288744101613345e+17, 1.288744101652407e+17, 1.288744101693033e+17, 1.288744101732096e+17, 1.288744101772719e+17, 1.288744101813345e+17, 1.288744101852407e+17, 1.288744101893032e+17, 1.288744101932095e+17, 1.288744101972719e+17, 1.288744102013345e+17, 1.288744102052407e+17, 1.288744102093033e+17, 1.288744102132095e+17, 1.288744102172719e+17, 1.288744102213345e+17, 1.288744102252407e+17, 1.288744102293033e+17, 1.288744102332095e+17, 1.288744102372719e+17, 1.288744102413345e+17, 1.288744102452407e+17, 1.288744102493033e+17, 1.288744102532095e+17, 1.288744102572721e+17, 1.288744102613345e+17, 1.288744102652407e+17, 1.288744102693033e+17, 1.288744102732095e+17, 1.288744102772719e+17, 1.288744102813345e+17, 1.288744102852407e+17, 1.288744102893033e+17, 1.288744102932095e+17, 1.288744102972721e+17, 1.288744103013345e+17, 1.288744103052407e+17, 1.288744103093033e+17, 1.288744103132095e+17, 1.288744103172721e+17, 1.288744103213345e+17, 1.288744103252407e+17, 1.288744103293033e+17, 1.288744103332095e+17, 1.288744103372721e+17, 1.288744103413344e+17, 1.288744103452408e+17, 1.288744103493033e+17, 1.288744103532095e+17, 1.288744103572721e+17, 1.288744103613344e+17, 1.288744103652407e+17, 1.288744103693032e+17, 1.288744103732095e+17, 1.288744103772721e+17, 1.288744103813345e+17, 1.288744103852408e+17, 1.288744103893032e+17, 1.288744103932096e+17, 1.288744103972719e+17, 1.288744104013344e+17, 1.288744104052408e+17, 1.288744104093032e+17, 1.288744104132095e+17, 1.288744104172719e+17, 1.288744104213345e+17, 1.288744104252407e+17, 1.288744104293033e+17, 1.288744104332096e+17, 1.288744104372719e+17, 1.288744104413345e+17, 1.288744104452407e+17, 1.288744104493032e+17, 1.288744104532095e+17, 1.288744104572719e+17, 1.288744104613345e+17, 1.288744104652407e+17, 1.288744104693033e+17, 1.288744104732095e+17, 1.288744104772719e+17, 1.288744104813345e+17, 1.288744104852407e+17, 1.288744104893033e+17, 1.288744104932095e+17, 1.288744104972719e+17, 1.288744105013345e+17, 1.288744105052407e+17, 1.288744105093033e+17, 1.288744105132095e+17, 1.288744105172721e+17, 1.288744105213345e+17, 1.288744105252407e+17, 1.288744105293033e+17, 1.288744105332095e+17, 1.288744105372719e+17, 1.288744105413345e+17, 1.288744105452407e+17, 1.288744105493033e+17, 1.288744105532095e+17, 1.288744105572721e+17, 1.288744105613345e+17, 1.288744105652408e+17, 1.288744105693033e+17, 1.288744105732095e+17, 1.288744105772721e+17, 1.288744105813345e+17, 1.288744105852407e+17, 1.288744105893033e+17, 1.288744105932095e+17, 1.288744105972721e+17, 1.288744106013345e+17, 1.288744106052408e+17, 1.288744106093033e+17, 1.288744106132095e+17, 1.288744106172721e+17, 1.288744106213344e+17, 1.288744106252407e+17, 1.288744106293032e+17, 1.288744106332095e+17, 1.288744106372721e+17, 1.288744106413345e+17, 1.288744106452408e+17, 1.288744106493032e+17, 1.288744106532096e+17, 1.288744106572719e+17, 1.288744106613345e+17, 1.288744106652408e+17, 1.288744106693032e+17, 1.288744106732095e+17, 1.288744106772719e+17, 1.288744106813345e+17, 1.288744106852407e+17, 1.288744106893033e+17, 1.288744106932096e+17, 1.288744106972719e+17, 1.288744107013345e+17, 1.288744107052407e+17, 1.288744107093032e+17, 1.288744107132095e+17, 1.288744107172719e+17, 1.288744107213345e+17, 1.288744107252407e+17, 1.288744107293033e+17, 1.288744107332095e+17, 1.288744107372719e+17, 1.288744107413345e+17, 1.288744107452407e+17, 1.288744107493033e+17, 1.288744107532095e+17, 1.288744107572719e+17, 1.288744107613345e+17, 1.288744107652407e+17, 1.288744107693033e+17, 1.288744107732095e+17, 1.288744107772721e+17, 1.288744107813345e+17, 1.288744107852407e+17, 1.288744107893033e+17, 1.288744107932095e+17, 1.288744107972719e+17, 1.288744108013345e+17, 1.288744108052407e+17, 1.288744108093033e+17, 1.288744108132095e+17, 1.288744108172721e+17, 1.288744108213345e+17, 1.288744108252408e+17, 1.288744108293033e+17, 1.288744108332095e+17, 1.288744108372721e+17, 1.288744108413344e+17, 1.288744108452407e+17, 1.288744108493033e+17, 1.288744108532095e+17, 1.288744108572721e+17, 1.288744108613345e+17, 1.288744108652408e+17, 1.288744108693032e+17, 1.288744108732095e+17, 1.288744108772721e+17, 1.288744108813344e+17, 1.288744108852408e+17, 1.288744108893032e+17, 1.288744108932095e+17, 1.288744108972719e+17, 1.288744109013345e+17, 1.288744109052408e+17, 1.288744109093032e+17, 1.288744109132096e+17, 1.288744109172719e+17, 1.288744109213345e+17, 1.288744109252407e+17, 1.288744109293032e+17, 1.288744109332095e+17, 1.288744109372719e+17, 1.288744109413345e+17, 1.288744109452407e+17, 1.288744109493033e+17, 1.288744109532095e+17, 1.288744109572719e+17, 1.288744109613345e+17, 1.288744109652407e+17, 1.288744109693032e+17, 1.288744109732095e+17, 1.288744109772719e+17, 1.288744109813345e+17, 1.288744109852407e+17, 1.288744109893033e+17, 1.288744109932095e+17, 1.288744109972719e+17, 1.288744110013345e+17, 1.288744110052407e+17, 1.288744110093033e+17, 1.288744110132095e+17, 1.288744110172719e+17, 1.288744110213345e+17, 1.288744110252407e+17, 1.288744110293033e+17, 1.288744110332095e+17, 1.288744110372721e+17, 1.288744110413345e+17, 1.288744110452407e+17, 1.288744110493033e+17, 1.288744110532095e+17, 1.288744110572719e+17, 1.288744110613345e+17, 1.288744110652407e+17, 1.288744110693033e+17, 1.288744110732095e+17, 1.288744110772721e+17, 1.288744110813345e+17, 1.288744110852408e+17, 1.288744110893033e+17, 1.288744110932095e+17, 1.288744110972721e+17, 1.288744111013344e+17, 1.288744111052407e+17, 1.288744111093033e+17, 1.288744111132095e+17, 1.288744111172721e+17, 1.288744111213345e+17, 1.288744111252408e+17, 1.288744111293032e+17, 1.288744111332095e+17, 1.288744111372721e+17, 1.288744111413344e+17, 1.288744111452408e+17, 1.288744111493032e+17, 1.288744111532095e+17, 1.288744111572719e+17, 1.288744111613345e+17, 1.288744111652408e+17, 1.288744111693032e+17, 1.288744111732096e+17, 1.288744111772719e+17, 1.288744111813345e+17, 1.288744111852407e+17, 1.288744111893032e+17, 1.288744111932095e+17, 1.288744111972719e+17, 1.288744112013345e+17, 1.288744112052407e+17, 1.288744112093033e+17, 1.288744112132095e+17, 1.288744112172719e+17, 1.288744112213345e+17, 1.288744112252407e+17, 1.288744112293032e+17, 1.288744112332095e+17, 1.288744112372719e+17, 1.288744112413345e+17, 1.288744112452407e+17, 1.288744112493033e+17, 1.288744112532095e+17, 1.288744112572721e+17, 1.288744112613345e+17, 1.288744112652407e+17, 1.288744112693033e+17, 1.288744112732095e+17, 1.288744112772719e+17, 1.288744112813345e+17, 1.288744112852407e+17, 1.288744112893033e+17, 1.288744112932095e+17, 1.288744112972721e+17, 1.288744113013345e+17, 1.288744113052407e+17, 1.288744113093033e+17, 1.288744113132095e+17, 1.288744113172719e+17, 1.288744113213345e+17, 1.288744113252407e+17, 1.288744113293033e+17, 1.288744113332095e+17, 1.288744113372721e+17, 1.288744113413345e+17, 1.288744113452408e+17, 1.288744113493033e+17, 1.288744113532095e+17, 1.288744113572721e+17, 1.288744113613344e+17, 1.288744113652407e+17, 1.288744113693033e+17, 1.288744113732095e+17, 1.288744113772721e+17, 1.288744113813345e+17, 1.288744113852408e+17, 1.288744113893032e+17, 1.288744113932095e+17, 1.288744113972721e+17, 1.288744114013344e+17, 1.288744114052408e+17, 1.288744114093032e+17, 1.288744114132095e+17, 1.288744114172719e+17, 1.288744114213345e+17, 1.288744114252408e+17, 1.288744114293032e+17, 1.288744114332096e+17, 1.288744114372719e+17, 1.288744114413345e+17, 1.288744114452407e+17, 1.288744114493032e+17, 1.288744114532095e+17, 1.288744114572719e+17, 1.288744114613345e+17, 1.288744114652407e+17, 1.288744114693033e+17, 1.288744114732095e+17, 1.288744114772719e+17, 1.288744114813345e+17, 1.288744114852407e+17, 1.288744114893032e+17, 1.288744114932095e+17, 1.288744114972719e+17, 1.288744115013345e+17, 1.288744115052407e+17, 1.288744115093033e+17, 1.288744115132095e+17, 1.288744115172721e+17, 1.288744115213345e+17, 1.288744115252407e+17, 1.288744115293033e+17, 1.288744115332095e+17, 1.288744115372719e+17, 1.288744115413345e+17, 1.288744115452407e+17, 1.288744115493033e+17, 1.288744115532095e+17, 1.288744115572721e+17, 1.288744115613345e+17, 1.288744115652407e+17, 1.288744115693033e+17, 1.288744115732095e+17, 1.288744115772721e+17, 1.288744115813345e+17, 1.288744115852407e+17, 1.288744115893033e+17, 1.288744115932095e+17, 1.288744115972721e+17, 1.288744116013344e+17, 1.288744116052408e+17, 1.288744116093033e+17, 1.288744116132095e+17, 1.288744116172721e+17, 1.288744116213344e+17, 1.288744116252407e+17, 1.288744116293032e+17, 1.288744116332095e+17, 1.288744116372721e+17, 1.288744116413345e+17, 1.288744116452408e+17, 1.288744116493032e+17, 1.288744116532095e+17, 1.288744116572719e+17, 1.288744116613344e+17, 1.288744116652408e+17, 1.288744116693032e+17, 1.288744116732095e+17, 1.288744116772719e+17, 1.288744116813345e+17, 1.288744116852407e+17, 1.288744116893032e+17, 1.288744116932096e+17, 1.288744116972719e+17, 1.288744117013345e+17, 1.288744117052407e+17, 1.288744117093032e+17, 1.288744117132095e+17, 1.288744117172719e+17, 1.288744117213345e+17, 1.288744117252407e+17, 1.288744117293033e+17, 1.288744117332095e+17, 1.288744117372719e+17, 1.288744117413345e+17, 1.288744117452407e+17, 1.288744117493032e+17, 1.288744117532095e+17, 1.288744117572719e+17, 1.288744117613345e+17, 1.288744117652407e+17, 1.288744117693033e+17, 1.288744117732095e+17, 1.288744117772721e+17, 1.288744117813345e+17, 1.288744117852407e+17, 1.288744117893033e+17, 1.288744117932095e+17, 1.288744117972719e+17, 1.288744118013345e+17, 1.288744118052407e+17, 1.288744118093033e+17, 1.288744118132095e+17, 1.288744118172721e+17, 1.288744118213345e+17, 1.288744118252407e+17, 1.288744118293033e+17, 1.288744118332095e+17, 1.288744118372721e+17, 1.288744118413345e+17, 1.288744118452407e+17, 1.288744118493033e+17, 1.288744118532095e+17, 1.288744118572721e+17, 1.288744118613344e+17, 1.288744118652408e+17, 1.288744118693033e+17, 1.288744118732095e+17, 1.288744118772721e+17, 1.288744118813344e+17, 1.288744118852407e+17, 1.288744118893032e+17, 1.288744118932095e+17, 1.288744118972721e+17, 1.288744119013345e+17, 1.288744119052408e+17, 1.288744119093032e+17, 1.288744119132096e+17, 1.288744119172719e+17, 1.288744119213344e+17, 1.288744119252408e+17, 1.288744119293032e+17, 1.288744119332095e+17, 1.288744119372719e+17, 1.288744119413345e+17, 1.288744119452407e+17, 1.288744119493033e+17, 1.288744119532096e+17, 1.288744119572719e+17, 1.288744119613345e+17, 1.288744119652407e+17, 1.288744119693032e+17, 1.288744119732095e+17, 1.288744119772719e+17, 1.288744119813345e+17, 1.288744119852407e+17, 1.288744119893033e+17, 1.288744119932095e+17, 1.288744119972719e+17, 1.288744120013345e+17, 1.288744120052407e+17, 1.288744120093033e+17, 1.288744120132095e+17, 1.288744120172719e+17, 1.288744120213345e+17, 1.288744120252407e+17, 1.288744120293033e+17, 1.288744120332095e+17, 1.288744120372721e+17, 1.288744120413345e+17, 1.288744120452407e+17, 1.288744120493033e+17, 1.288744120532095e+17, 1.288744120572719e+17, 1.288744120613345e+17, 1.288744120652407e+17, 1.288744120693033e+17, 1.288744120732095e+17, 1.288744120772721e+17, 1.288744120813345e+17, 1.288744120852407e+17, 1.288744120893033e+17, 1.288744120932095e+17, 1.288744120972721e+17, 1.288744121013345e+17, 1.288744121052407e+17, 1.288744121093033e+17, 1.288744121132095e+17, 1.288744121172721e+17, 1.288744121213344e+17, 1.288744121252408e+17, 1.288744121293033e+17, 1.288744121332095e+17, 1.288744121372721e+17, 1.288744121413344e+17, 1.288744121452407e+17, 1.288744121493032e+17, 1.288744121532095e+17, 1.288744121572721e+17, 1.288744121613345e+17, 1.288744121652408e+17, 1.288744121693032e+17, 1.288744121732096e+17, 1.288744121772719e+17, 1.288744121813344e+17, 1.288744121852408e+17, 1.288744121893032e+17, 1.288744121932095e+17, 1.288744121972719e+17, 1.288744122013345e+17, 1.288744122052407e+17, 1.288744122093033e+17, 1.288744122132096e+17, 1.288744122172719e+17, 1.288744122213345e+17, 1.288744122252407e+17, 1.288744122293032e+17, 1.288744122332095e+17, 1.288744122372719e+17, 1.288744122413345e+17, 1.288744122452407e+17, 1.288744122493033e+17, 1.288744122532095e+17, 1.288744122572719e+17, 1.288744122613345e+17, 1.288744122652407e+17, 1.288744122693033e+17, 1.288744122732095e+17, 1.288744122772719e+17, 1.288744122813345e+17, 1.288744122852407e+17, 1.288744122893033e+17, 1.288744122932095e+17, 1.288744122972721e+17, 1.288744123013345e+17, 1.288744123052407e+17, 1.288744123093033e+17, 1.288744123132095e+17, 1.288744123172719e+17, 1.288744123213345e+17, 1.288744123252407e+17, 1.288744123293033e+17, 1.288744123332095e+17, 1.288744123372721e+17, 1.288744123413345e+17, 1.288744123452407e+17, 1.288744123493033e+17, 1.288744123532095e+17, 1.288744123572721e+17, 1.288744123613345e+17, 1.288744123652407e+17, 1.288744123693033e+17, 1.288744123732095e+17, 1.288744123772721e+17, 1.288744123813345e+17, 1.288744123852408e+17, 1.288744123893033e+17, 1.288744123932095e+17, 1.288744123972721e+17, 1.288744124013344e+17, 1.288744124052407e+17, 1.288744124093032e+17, 1.288744124132095e+17, 1.288744124172721e+17, 1.288744124213345e+17, 1.288744124252408e+17, 1.288744124293032e+17, 1.288744124332096e+17, 1.288744124372719e+17, 1.288744124413344e+17, 1.288744124452408e+17, 1.288744124493032e+17, 1.288744124532095e+17, 1.288744124572719e+17, 1.288744124613345e+17, 1.288744124652407e+17, 1.288744124693033e+17, 1.288744124732096e+17, 1.288744124772719e+17, 1.288744124813345e+17, 1.288744124852407e+17, 1.288744124893032e+17, 1.288744124932095e+17, 1.288744124972719e+17, 1.288744125013345e+17, 1.288744125052407e+17, 1.288744125093033e+17, 1.288744125132095e+17, 1.288744125172719e+17, 1.288744125213345e+17, 1.288744125252407e+17, 1.288744125293033e+17, 1.288744125332095e+17, 1.288744125372719e+17, 1.288744125413345e+17, 1.288744125452407e+17, 1.288744125493033e+17, 1.288744125532095e+17, 1.288744125572721e+17, 1.288744125613345e+17, 1.288744125652407e+17, 1.288744125693033e+17, 1.288744125732095e+17, 1.288744125772719e+17, 1.288744125813345e+17, 1.288744125852407e+17, 1.288744125893033e+17, 1.288744125932095e+17, 1.288744125972721e+17, 1.288744126013345e+17, 1.288744126052408e+17, 1.288744126093033e+17, 1.288744126132095e+17, 1.288744126172721e+17, 1.288744126213344e+17, 1.288744126252407e+17, 1.288744126293033e+17, 1.288744126332095e+17, 1.288744126372721e+17, 1.288744126413345e+17, 1.288744126452408e+17, 1.288744126493032e+17, 1.288744126532095e+17, 1.288744126572721e+17, 1.288744126613344e+17, 1.288744126652408e+17, 1.288744126693032e+17, 1.288744126732095e+17, 1.288744126772719e+17, 1.288744126813345e+17, 1.288744126852408e+17, 1.288744126893032e+17, 1.288744126932096e+17, 1.288744126972719e+17, 1.288744127013345e+17, 1.288744127052407e+17, 1.288744127093032e+17, 1.288744127132095e+17, 1.288744127172719e+17, 1.288744127213345e+17, 1.288744127252407e+17, 1.288744127293033e+17, 1.288744127332095e+17, 1.288744127372719e+17, 1.288744127413345e+17, 1.288744127452407e+17, 1.288744127493032e+17, 1.288744127532095e+17, 1.288744127572719e+17, 1.288744127613345e+17, 1.288744127652407e+17, 1.288744127693033e+17, 1.288744127732095e+17, 1.288744127772719e+17, 1.288744127813345e+17, 1.288744127852407e+17, 1.288744127893033e+17, 1.288744127932095e+17, 1.288744127972719e+17, 1.288744128013345e+17, 1.288744128052407e+17, 1.288744128093033e+17, 1.288744128132095e+17, 1.288744128172721e+17, 1.288744128213345e+17, 1.288744128252407e+17, 1.288744128293033e+17, 1.288744128332095e+17, 1.288744128372719e+17, 1.288744128413345e+17, 1.288744128452407e+17, 1.288744128493033e+17, 1.288744128532095e+17, 1.288744128572721e+17, 1.288744128613345e+17, 1.288744128652408e+17, 1.288744128693033e+17, 1.288744128732095e+17, 1.288744128772721e+17, 1.288744128813344e+17, 1.288744128852407e+17, 1.288744128893033e+17, 1.288744128932095e+17, 1.288744128972721e+17, 1.288744129013345e+17, 1.288744129052408e+17, 1.288744129093032e+17, 1.288744129132095e+17, 1.288744129172721e+17, 1.288744129213344e+17, 1.288744129252408e+17, 1.288744129293032e+17, 1.288744129332095e+17, 1.288744129372719e+17, 1.288744129413345e+17, 1.288744129452408e+17, 1.288744129493032e+17, 1.288744129532096e+17, 1.288744129572719e+17, 1.288744129613345e+17, 1.288744129652407e+17, 1.288744129693032e+17, 1.288744129732095e+17, 1.288744129772719e+17, 1.288744129813345e+17, 1.288744129852407e+17, 1.288744129893033e+17, 1.288744129932095e+17, 1.288744129972719e+17, 1.288744130013345e+17, 1.288744130052407e+17, 1.288744130093032e+17, 1.288744130132095e+17, 1.288744130172719e+17, 1.288744130213345e+17, 1.288744130252407e+17, 1.288744130293033e+17, 1.288744130332095e+17, 1.288744130372719e+17, 1.288744130413345e+17, 1.288744130452407e+17, 1.288744130493033e+17, 1.288744130532095e+17, 1.288744130572719e+17, 1.288744130613345e+17, 1.288744130652407e+17, 1.288744130693033e+17, 1.288744130732095e+17, 1.288744130772721e+17, 1.288744130813345e+17, 1.288744130852407e+17, 1.288744130893033e+17, 1.288744130932095e+17, 1.288744130972719e+17, 1.288744131013345e+17, 1.288744131052407e+17, 1.288744131093033e+17, 1.288744131132095e+17, 1.288744131172721e+17, 1.288744131213345e+17, 1.288744131252408e+17, 1.288744131293033e+17, 1.288744131332095e+17, 1.288744131372721e+17, 1.288744131413344e+17, 1.288744131452407e+17, 1.288744131493033e+17, 1.288744131532095e+17, 1.288744131572721e+17, 1.288744131613345e+17, 1.288744131652408e+17, 1.288744131693032e+17, 1.288744131732095e+17, 1.288744131772721e+17, 1.288744131813344e+17, 1.288744131852408e+17, 1.288744131893032e+17, 1.288744131932095e+17, 1.288744131972719e+17, 1.288744132013345e+17, 1.288744132052408e+17, 1.288744132093032e+17, 1.288744132132096e+17, 1.288744132172719e+17, 1.288744132213345e+17, 1.288744132252407e+17, 1.288744132293032e+17, 1.288744132332095e+17, 1.288744132372719e+17, 1.288744132413345e+17, 1.288744132452407e+17, 1.288744132493033e+17, 1.288744132532095e+17, 1.288744132572719e+17, 1.288744132613345e+17, 1.288744132652407e+17, 1.288744132693032e+17, 1.288744132732095e+17, 1.288744132772719e+17, 1.288744132813345e+17, 1.288744132852407e+17, 1.288744132893033e+17, 1.288744132932095e+17, 1.288744132972721e+17, 1.288744133013345e+17, 1.288744133052407e+17, 1.288744133093033e+17, 1.288744133132095e+17, 1.288744133172719e+17, 1.288744133213345e+17, 1.288744133252407e+17, 1.288744133293033e+17, 1.288744133332095e+17, 1.288744133372721e+17, 1.288744133413345e+17, 1.288744133452407e+17, 1.288744133493033e+17, 1.288744133532095e+17, 1.288744133572721e+17, 1.288744133613345e+17, 1.288744133652407e+17, 1.288744133693033e+17, 1.288744133732095e+17, 1.288744133772721e+17, 1.288744133813345e+17, 1.288744133852408e+17, 1.288744133893033e+17, 1.288744133932095e+17, 1.288744133972721e+17, 1.288744134013344e+17, 1.288744134052407e+17, 1.288744134093033e+17, 1.288744134132095e+17, 1.288744134172721e+17, 1.288744134213345e+17, 1.288744134252408e+17, 1.288744134293032e+17, 1.288744134332095e+17, 1.288744134372721e+17, 1.288744134413344e+17, 1.288744134452408e+17, 1.288744134493032e+17, 1.288744134532095e+17, 1.288744134572719e+17, 1.288744134613345e+17, 1.288744134652408e+17, 1.288744134693032e+17, 1.288744134732096e+17, 1.288744134772719e+17, 1.288744134813345e+17, 1.288744134852407e+17, 1.288744134893032e+17, 1.288744134932095e+17, 1.288744134972719e+17, 1.288744135013345e+17, 1.288744135052407e+17, 1.288744135093033e+17, 1.288744135132095e+17, 1.288744135172719e+17, 1.288744135213345e+17, 1.288744135252407e+17, 1.288744135293032e+17, 1.288744135332095e+17, 1.288744135372719e+17, 1.288744135413345e+17, 1.288744135452407e+17, 1.288744135493033e+17, 1.288744135532095e+17, 1.288744135572721e+17, 1.288744135613345e+17, 1.288744135652407e+17, 1.288744135693033e+17, 1.288744135732095e+17, 1.288744135772719e+17, 1.288744135813345e+17, 1.288744135852407e+17, 1.288744135893033e+17, 1.288744135932095e+17, 1.288744135972721e+17, 1.288744136013345e+17, 1.288744136052407e+17, 1.288744136093033e+17, 1.288744136132095e+17, 1.288744136172721e+17, 1.288744136213345e+17, 1.288744136252407e+17, 1.288744136293033e+17, 1.288744136332095e+17, 1.288744136372721e+17, 1.288744136413344e+17, 1.288744136452408e+17, 1.288744136493033e+17, 1.288744136532095e+17, 1.288744136572721e+17, 1.288744136613344e+17, 1.288744136652407e+17, 1.288744136693032e+17, 1.288744136732095e+17, 1.288744136772721e+17, 1.288744136813345e+17, 1.288744136852408e+17, 1.288744136893032e+17, 1.288744136932095e+17, 1.288744136972719e+17, 1.288744137013344e+17, 1.288744137052408e+17, 1.288744137093032e+17, 1.288744137132095e+17, 1.288744137172719e+17, 1.288744137213345e+17, 1.288744137252407e+17, 1.288744137293033e+17, 1.288744137332096e+17, 1.288744137372719e+17, 1.288744137413345e+17, 1.288744137452407e+17, 1.288744137493032e+17, 1.288744137532095e+17, 1.288744137572719e+17, 1.288744137613345e+17, 1.288744137652407e+17, 1.288744137693033e+17, 1.288744137732095e+17, 1.288744137772719e+17, 1.288744137813345e+17, 1.288744137852407e+17, 1.288744137893032e+17, 1.288744137932095e+17, 1.288744137972719e+17, 1.288744138013345e+17, 1.288744138052407e+17, 1.288744138093033e+17, 1.288744138132095e+17, 1.288744138172721e+17, 1.288744138213345e+17, 1.288744138252407e+17, 1.288744138293033e+17, 1.288744138332095e+17, 1.288744138372719e+17, 1.288744138413345e+17, 1.288744138452407e+17, 1.288744138493033e+17, 1.288744138532095e+17, 1.288744138572721e+17, 1.288744138613345e+17, 1.288744138652407e+17, 1.288744138693033e+17, 1.288744138732095e+17, 1.288744138772721e+17, 1.288744138813345e+17, 1.288744138852407e+17, 1.288744138893033e+17, 1.288744138932095e+17, 1.288744138972721e+17, 1.288744139013344e+17, 1.288744139052408e+17, 1.288744139093033e+17, 1.288744139132095e+17, 1.288744139172721e+17, 1.288744139213344e+17, 1.288744139252407e+17, 1.288744139293032e+17, 1.288744139332095e+17, 1.288744139372721e+17, 1.288744139413345e+17, 1.288744139452408e+17, 1.288744139493032e+17, 1.288744139532096e+17, 1.288744139572719e+17, 1.288744139613344e+17, 1.288744139652408e+17, 1.288744139693032e+17, 1.288744139732095e+17, 1.288744139772719e+17, 1.288744139813345e+17, 1.288744139852407e+17, 1.288744139893033e+17, 1.288744139932096e+17, 1.288744139972719e+17, 1.288744140013345e+17, 1.288744140052407e+17, 1.288744140093032e+17, 1.288744140132095e+17, 1.288744140172719e+17, 1.288744140213345e+17, 1.288744140252407e+17, 1.288744140293033e+17, 1.288744140332095e+17, 1.288744140372719e+17, 1.288744140413345e+17, 1.288744140452407e+17, 1.288744140493033e+17, 1.288744140532095e+17, 1.288744140572719e+17, 1.288744140613345e+17, 1.288744140652407e+17, 1.288744140693033e+17, 1.288744140732095e+17, 1.288744140772721e+17, 1.288744140813345e+17, 1.288744140852407e+17, 1.288744140893033e+17, 1.288744140932095e+17, 1.288744140972719e+17, 1.288744141013345e+17, 1.288744141052407e+17, 1.288744141093033e+17, 1.288744141132095e+17, 1.288744141172721e+17, 1.288744141213345e+17, 1.288744141252407e+17, 1.288744141293033e+17, 1.288744141332095e+17, 1.288744141372721e+17, 1.288744141413345e+17, 1.288744141452407e+17, 1.288744141493033e+17, 1.288744141532095e+17, 1.288744141572721e+17, 1.288744141613344e+17, 1.288744141652408e+17, 1.288744141693033e+17, 1.288744141732095e+17, 1.288744141772721e+17, 1.288744141813344e+17, 1.288744141852407e+17, 1.288744141893032e+17, 1.288744141932095e+17, 1.288744141972721e+17, 1.288744142013345e+17, 1.288744142052408e+17, 1.288744142093032e+17, 1.288744142132096e+17, 1.288744142172719e+17, 1.288744142213344e+17, 1.288744142252408e+17, 1.288744142293032e+17, 1.288744142332095e+17, 1.288744142372719e+17, 1.288744142413345e+17, 1.288744142452407e+17, 1.288744142493033e+17, 1.288744142532096e+17, 1.288744142572719e+17, 1.288744142613345e+17, 1.288744142652407e+17, 1.288744142693032e+17, 1.288744142732095e+17, 1.288744142772719e+17, 1.288744142813345e+17, 1.288744142852407e+17, 1.288744142893033e+17, 1.288744142932095e+17, 1.288744142972719e+17, 1.288744143013345e+17, 1.288744143052407e+17, 1.288744143093033e+17, 1.288744143132095e+17, 1.288744143172719e+17, 1.288744143213345e+17, 1.288744143252407e+17, 1.288744143293033e+17, 1.288744143332095e+17, 1.288744143372721e+17, 1.288744143413345e+17, 1.288744143452407e+17, 1.288744143493033e+17, 1.288744143532095e+17, 1.288744143572719e+17, 1.288744143613345e+17, 1.288744143652407e+17, 1.288744143693033e+17, 1.288744143732095e+17, 1.288744143772721e+17, 1.288744143813345e+17, 1.288744143852408e+17, 1.288744143893033e+17, 1.288744143932095e+17, 1.288744143972721e+17, 1.288744144013345e+17, 1.288744144052407e+17, 1.288744144093033e+17, 1.288744144132095e+17, 1.288744144172721e+17, 1.288744144213345e+17, 1.288744144252408e+17, 1.288744144293033e+17, 1.288744144332095e+17, 1.288744144372721e+17, 1.288744144413344e+17, 1.288744144452407e+17, 1.288744144493032e+17, 1.288744144532095e+17, 1.288744144572721e+17, 1.288744144613345e+17, 1.288744144652408e+17, 1.288744144693032e+17, 1.288744144732096e+17, 1.288744144772719e+17, 1.288744144813344e+17, 1.288744144852408e+17, 1.288744144893032e+17, 1.288744144932095e+17, 1.288744144972719e+17, 1.288744145013345e+17, 1.288744145052407e+17, 1.288744145093033e+17, 1.288744145132096e+17, 1.288744145172719e+17, 1.288744145213345e+17, 1.288744145252407e+17, 1.288744145293032e+17, 1.288744145332095e+17, 1.288744145372719e+17, 1.288744145413345e+17, 1.288744145452407e+17, 1.288744145493033e+17, 1.288744145532095e+17, 1.288744145572719e+17, 1.288744145613345e+17, 1.288744145652407e+17, 1.288744145693033e+17, 1.288744145732095e+17, 1.288744145772719e+17, 1.288744145813345e+17, 1.288744145852407e+17, 1.288744145893033e+17, 1.288744145932095e+17, 1.288744145972721e+17, 1.288744146013345e+17, 1.288744146052407e+17, 1.288744146093033e+17, 1.288744146132095e+17, 1.288744146172719e+17, 1.288744146213345e+17, 1.288744146252407e+17, 1.288744146293033e+17, 1.288744146332095e+17, 1.288744146372721e+17, 1.288744146413345e+17, 1.288744146452408e+17, 1.288744146493033e+17, 1.288744146532095e+17, 1.288744146572721e+17, 1.288744146613344e+17, 1.288744146652407e+17, 1.288744146693033e+17, 1.288744146732095e+17, 1.288744146772721e+17, 1.288744146813345e+17, 1.288744146852408e+17, 1.288744146893032e+17, 1.288744146932095e+17, 1.288744146972721e+17, 1.288744147013344e+17, 1.288744147052408e+17, 1.288744147093032e+17, 1.288744147132095e+17, 1.288744147172719e+17, 1.288744147213345e+17, 1.288744147252408e+17, 1.288744147293032e+17, 1.288744147332096e+17, 1.288744147372719e+17, 1.288744147413345e+17, 1.288744147452407e+17, 1.288744147493032e+17, 1.288744147532095e+17, 1.288744147572719e+17, 1.288744147613345e+17, 1.288744147652407e+17, 1.288744147693033e+17, 1.288744147732095e+17, 1.288744147772719e+17, 1.288744147813345e+17, 1.288744147852407e+17, 1.288744147893032e+17, 1.288744147932095e+17, 1.288744147972719e+17, 1.288744148013345e+17, 1.288744148052407e+17, 1.288744148093033e+17, 1.288744148132095e+17, 1.288744148172719e+17, 1.288744148213345e+17, 1.288744148252407e+17, 1.288744148293033e+17, 1.288744148332095e+17, 1.288744148372719e+17, 1.288744148413345e+17, 1.288744148452407e+17, 1.288744148493033e+17, 1.288744148532095e+17, 1.288744148572721e+17, 1.288744148613345e+17, 1.288744148652407e+17, 1.288744148693033e+17, 1.288744148732095e+17, 1.288744148772719e+17, 1.288744148813345e+17, 1.288744148852407e+17, 1.288744148893033e+17, 1.288744148932095e+17, 1.288744148972721e+17, 1.288744149013345e+17, 1.288744149052408e+17, 1.288744149093033e+17, 1.288744149132095e+17, 1.288744149172721e+17, 1.288744149213344e+17, 1.288744149252407e+17, 1.288744149293033e+17, 1.288744149332095e+17, 1.288744149372721e+17, 1.288744149413345e+17, 1.288744149452408e+17, 1.288744149493032e+17, 1.288744149532095e+17, 1.288744149572721e+17, 1.288744149613344e+17, 1.288744149652408e+17, 1.288744149693032e+17, 1.288744149732095e+17, 1.288744149772719e+17, 1.288744149813345e+17, 1.288744149852408e+17, 1.288744149893032e+17, 1.288744149932096e+17, 1.288744149972719e+17, 1.288744150013345e+17, 1.288744150052407e+17, 1.288744150093032e+17, 1.288744150132095e+17, 1.288744150172719e+17, 1.288744150213345e+17, 1.288744150252407e+17, 1.288744150293033e+17, 1.288744150332095e+17, 1.288744150372719e+17, 1.288744150413345e+17, 1.288744150452407e+17, 1.288744150493032e+17, 1.288744150532095e+17, 1.288744150572719e+17, 1.288744150613345e+17, 1.288744150652407e+17, 1.288744150693033e+17, 1.288744150732095e+17, 1.288744150772721e+17, 1.288744150813345e+17, 1.288744150852407e+17, 1.288744150893033e+17, 1.288744150932095e+17, 1.288744150972719e+17, 1.288744151013345e+17, 1.288744151052407e+17, 1.288744151093033e+17, 1.288744151132095e+17, 1.288744151172721e+17, 1.288744151213345e+17, 1.288744151252407e+17, 1.288744151293033e+17, 1.288744151332095e+17, 1.288744151372719e+17, 1.288744151413345e+17, 1.288744151452407e+17, 1.288744151493033e+17, 1.288744151532095e+17, 1.288744151572721e+17, 1.288744151613345e+17, 1.288744151652408e+17, 1.288744151693033e+17, 1.288744151732095e+17, 1.288744151772721e+17, 1.288744151813344e+17, 1.288744151852407e+17, 1.288744151893033e+17, 1.288744151932095e+17, 1.288744151972721e+17, 1.288744152013345e+17, 1.288744152052408e+17, 1.288744152093032e+17, 1.288744152132095e+17, 1.288744152172721e+17, 1.288744152213344e+17, 1.288744152252408e+17, 1.288744152293032e+17, 1.288744152332095e+17, 1.288744152372719e+17, 1.288744152413345e+17, 1.288744152452408e+17, 1.288744152493032e+17, 1.288744152532096e+17, 1.288744152572719e+17, 1.288744152613345e+17, 1.288744152652407e+17, 1.288744152693032e+17, 1.288744152732095e+17, 1.288744152772719e+17, 1.288744152813345e+17, 1.288744152852407e+17, 1.288744152893033e+17, 1.288744152932095e+17, 1.288744152972719e+17, 1.288744153013345e+17, 1.288744153052407e+17, 1.288744153093032e+17, 1.288744153132095e+17, 1.288744153172719e+17, 1.288744153213345e+17, 1.288744153252407e+17, 1.288744153293033e+17, 1.288744153332095e+17, 1.288744153372721e+17, 1.288744153413345e+17, 1.288744153452407e+17, 1.288744153493033e+17, 1.288744153532095e+17, 1.288744153572719e+17, 1.288744153613345e+17, 1.288744153652407e+17, 1.288744153693033e+17, 1.288744153732095e+17, 1.288744153772721e+17, 1.288744153813345e+17, 1.288744153852407e+17, 1.288744153893033e+17, 1.288744153932095e+17, 1.288744153972721e+17, 1.288744154013345e+17, 1.288744154052407e+17, 1.288744154093033e+17, 1.288744154132095e+17, 1.288744154172721e+17, 1.288744154213345e+17, 1.288744154252408e+17, 1.288744154293033e+17, 1.288744154332095e+17, 1.288744154372721e+17, 1.288744154413344e+17, 1.288744154452407e+17, 1.288744154493033e+17, 1.288744154532095e+17, 1.288744154572721e+17, 1.288744154613345e+17, 1.288744154652408e+17, 1.288744154693032e+17, 1.288744154732095e+17, 1.288744154772721e+17, 1.288744154813344e+17, 1.288744154852408e+17, 1.288744154893032e+17, 1.288744154932095e+17, 1.288744154972719e+17, 1.288744155013345e+17, 1.288744155052408e+17, 1.288744155093032e+17, 1.288744155132096e+17, 1.288744155172719e+17, 1.288744155213345e+17, 1.288744155252407e+17, 1.288744155293032e+17, 1.288744155332095e+17, 1.288744155372719e+17, 1.288744155413345e+17, 1.288744155452407e+17, 1.288744155493033e+17, 1.288744155532095e+17, 1.288744155572719e+17, 1.288744155613345e+17, 1.288744155652407e+17, 1.288744155693032e+17, 1.288744155732095e+17, 1.288744155772719e+17, 1.288744155813345e+17, 1.288744155852407e+17, 1.288744155893033e+17, 1.288744155932095e+17, 1.288744155972721e+17, 1.288744156013345e+17, 1.288744156052407e+17, 1.288744156093033e+17, 1.288744156132095e+17, 1.288744156172719e+17, 1.288744156213345e+17, 1.288744156252407e+17, 1.288744156293033e+17, 1.288744156332095e+17, 1.288744156372721e+17, 1.288744156413345e+17, 1.288744156452407e+17, 1.288744156493033e+17, 1.288744156532095e+17, 1.288744156572721e+17, 1.288744156613345e+17, 1.288744156652407e+17, 1.288744156693033e+17, 1.288744156732095e+17, 1.288744156772721e+17, 1.288744156813344e+17, 1.288744156852408e+17, 1.288744156893033e+17, 1.288744156932095e+17, 1.288744156972721e+17, 1.288744157013344e+17, 1.288744157052407e+17, 1.288744157093032e+17, 1.288744157132095e+17, 1.288744157172721e+17, 1.288744157213345e+17, 1.288744157252408e+17, 1.288744157293032e+17, 1.288744157332096e+17, 1.288744157372719e+17, 1.288744157413344e+17, 1.288744157452408e+17, 1.288744157493032e+17, 1.288744157532095e+17, 1.288744157572719e+17, 1.288744157613345e+17, 1.288744157652407e+17, 1.288744157693033e+17, 1.288744157732096e+17, 1.288744157772719e+17, 1.288744157813345e+17, 1.288744157852407e+17, 1.288744157893032e+17, 1.288744157932095e+17, 1.288744157972719e+17, 1.288744158013345e+17, 1.288744158052407e+17, 1.288744158093033e+17, 1.288744158132095e+17, 1.288744158172719e+17, 1.288744158213345e+17, 1.288744158252407e+17, 1.288744158293033e+17, 1.288744158332095e+17, 1.288744158372719e+17, 1.288744158413345e+17, 1.288744158452407e+17, 1.288744158493033e+17, 1.288744158532095e+17, 1.288744158572721e+17, 1.288744158613345e+17, 1.288744158652407e+17, 1.288744158693033e+17, 1.288744158732095e+17, 1.288744158772719e+17, 1.288744158813345e+17, 1.288744158852407e+17, 1.288744158893033e+17, 1.288744158932095e+17, 1.288744158972721e+17, 1.288744159013345e+17, 1.288744159052407e+17, 1.288744159093033e+17, 1.288744159132095e+17, 1.288744159172721e+17, 1.288744159213345e+17, 1.288744159252407e+17, 1.288744159293033e+17, 1.288744159332095e+17, 1.288744159372721e+17, 1.288744159413344e+17, 1.288744159452408e+17, 1.288744159493033e+17, 1.288744159532095e+17, 1.288744159572721e+17, 1.288744159613344e+17, 1.288744159652407e+17, 1.288744159693032e+17, 1.288744159732095e+17, 1.288744159772721e+17, 1.288744159813345e+17, 1.288744159852408e+17, 1.288744159893032e+17, 1.288744159932096e+17, 1.288744159972719e+17, 1.288744160013344e+17, 1.288744160052408e+17, 1.288744160093032e+17, 1.288744160132095e+17, 1.288744160172719e+17, 1.288744160213345e+17, 1.288744160252407e+17, 1.288744160293033e+17, 1.288744160332096e+17, 1.288744160372719e+17, 1.288744160413345e+17, 1.288744160452407e+17, 1.288744160493032e+17, 1.288744160532095e+17, 1.288744160572719e+17, 1.288744160613345e+17, 1.288744160652407e+17, 1.288744160693033e+17, 1.288744160732095e+17, 1.288744160772719e+17, 1.288744160813345e+17, 1.288744160852407e+17, 1.288744160893033e+17, 1.288744160932095e+17, 1.288744160972719e+17, 1.288744161013345e+17, 1.288744161052407e+17, 1.288744161093033e+17, 1.288744161132095e+17, 1.288744161172721e+17, 1.288744161213345e+17, 1.288744161252407e+17, 1.288744161293033e+17, 1.288744161332095e+17, 1.288744161372719e+17, 1.288744161413345e+17, 1.288744161452407e+17, 1.288744161493033e+17, 1.288744161532095e+17, 1.288744161572721e+17, 1.288744161613345e+17, 1.288744161652407e+17, 1.288744161693033e+17, 1.288744161732095e+17, 1.288744161772721e+17, 1.288744161813345e+17, 1.288744161852407e+17, 1.288744161893033e+17, 1.288744161932095e+17, 1.288744161972721e+17, 1.288744162013344e+17, 1.288744162052408e+17, 1.288744162093033e+17, 1.288744162132095e+17, 1.288744162172721e+17, 1.288744162213344e+17, 1.288744162252407e+17, 1.288744162293032e+17, 1.288744162332095e+17, 1.288744162372721e+17, 1.288744162413345e+17, 1.288744162452408e+17, 1.288744162493032e+17, 1.288744162532096e+17, 1.288744162572719e+17, 1.288744162613344e+17, 1.288744162652408e+17, 1.288744162693032e+17, 1.288744162732095e+17, 1.288744162772719e+17, 1.288744162813345e+17, 1.288744162852407e+17, 1.288744162893033e+17, 1.288744162932096e+17, 1.288744162972719e+17, 1.288744163013345e+17, 1.288744163052407e+17, 1.288744163093032e+17, 1.288744163132095e+17, 1.288744163172719e+17, 1.288744163213345e+17, 1.288744163252407e+17, 1.288744163293033e+17, 1.288744163332095e+17, 1.288744163372719e+17, 1.288744163413345e+17, 1.288744163452407e+17, 1.288744163493033e+17, 1.288744163532095e+17, 1.288744163572719e+17, 1.288744163613345e+17, 1.288744163652407e+17, 1.288744163693033e+17, 1.288744163732095e+17, 1.288744163772721e+17, 1.288744163813345e+17, 1.288744163852407e+17, 1.288744163893033e+17, 1.288744163932095e+17, 1.288744163972719e+17, 1.288744164013345e+17, 1.288744164052407e+17, 1.288744164093033e+17, 1.288744164132095e+17, 1.288744164172721e+17, 1.288744164213345e+17, 1.288744164252408e+17, 1.288744164293033e+17, 1.288744164332095e+17, 1.288744164372721e+17, 1.288744164413344e+17, 1.288744164452407e+17, 1.288744164493033e+17, 1.288744164532095e+17, 1.288744164572721e+17, 1.288744164613345e+17, 1.288744164652408e+17, 1.288744164693032e+17, 1.288744164732095e+17, 1.288744164772721e+17, 1.288744164813344e+17, 1.288744164852407e+17, 1.288744164893032e+17, 1.288744164932095e+17, 1.288744164972719e+17, 1.288744165013345e+17, 1.288744165052408e+17, 1.288744165093032e+17, 1.288744165132096e+17, 1.288744165172719e+17, 1.288744165213345e+17, 1.288744165252407e+17, 1.288744165293032e+17, 1.288744165332095e+17, 1.288744165372719e+17, 1.288744165413345e+17, 1.288744165452407e+17, 1.288744165493033e+17, 1.288744165532095e+17, 1.288744165572719e+17, 1.288744165613345e+17, 1.288744165652407e+17, 1.288744165693032e+17, 1.288744165732095e+17, 1.288744165772719e+17, 1.288744165813345e+17, 1.288744165852407e+17, 1.288744165893033e+17, 1.288744165932095e+17, 1.288744165972719e+17, 1.288744166013345e+17, 1.288744166052407e+17, 1.288744166093033e+17, 1.288744166132095e+17, 1.288744166172719e+17, 1.288744166213345e+17, 1.288744166252407e+17, 1.288744166293033e+17, 1.288744166332095e+17, 1.288744166372721e+17, 1.288744166413345e+17, 1.288744166452407e+17, 1.288744166493033e+17, 1.288744166532095e+17, 1.288744166572719e+17, 1.288744166613345e+17, 1.288744166652407e+17, 1.288744166693033e+17, 1.288744166732095e+17, 1.288744166772721e+17, 1.288744166813345e+17, 1.288744166852408e+17, 1.288744166893033e+17, 1.288744166932095e+17, 1.288744166972721e+17, 1.288744167013344e+17, 1.288744167052407e+17, 1.288744167093033e+17, 1.288744167132095e+17, 1.288744167172721e+17, 1.288744167213345e+17, 1.288744167252408e+17, 1.288744167293032e+17, 1.288744167332095e+17, 1.288744167372721e+17, 1.288744167413344e+17, 1.288744167452408e+17, 1.288744167493032e+17, 1.288744167532095e+17, 1.288744167572719e+17, 1.288744167613345e+17, 1.288744167652408e+17, 1.288744167693032e+17, 1.288744167732096e+17, 1.288744167772719e+17, 1.288744167813345e+17, 1.288744167852407e+17, 1.288744167893032e+17, 1.288744167932095e+17, 1.288744167972719e+17, 1.288744168013345e+17, 1.288744168052407e+17, 1.288744168093033e+17, 1.288744168132095e+17, 1.288744168172719e+17, 1.288744168213345e+17, 1.288744168252407e+17, 1.288744168293032e+17, 1.288744168332095e+17, 1.288744168372719e+17, 1.288744168413345e+17, 1.288744168452407e+17, 1.288744168493033e+17, 1.288744168532095e+17, 1.288744168572719e+17, 1.288744168613345e+17, 1.288744168652407e+17, 1.288744168693033e+17, 1.288744168732095e+17, 1.288744168772719e+17, 1.288744168813345e+17, 1.288744168852407e+17, 1.288744168893033e+17, 1.288744168932095e+17, 1.288744168972721e+17, 1.288744169013345e+17, 1.288744169052407e+17, 1.288744169093033e+17, 1.288744169132095e+17, 1.288744169172719e+17, 1.288744169213345e+17, 1.288744169252407e+17, 1.288744169293033e+17, 1.288744169332095e+17, 1.288744169372721e+17, 1.288744169413345e+17, 1.288744169452408e+17, 1.288744169493033e+17, 1.288744169532095e+17, 1.288744169572721e+17, 1.288744169613344e+17, 1.288744169652407e+17, 1.288744169693033e+17, 1.288744169732095e+17, 1.288744169772721e+17, 1.288744169813345e+17, 1.288744169852408e+17, 1.288744169893032e+17, 1.288744169932095e+17, 1.288744169972721e+17, 1.288744170013344e+17, 1.288744170052408e+17, 1.288744170093032e+17, 1.288744170132095e+17, 1.288744170172719e+17, 1.288744170213345e+17, 1.288744170252408e+17, 1.288744170293032e+17, 1.288744170332096e+17, 1.288744170372719e+17, 1.288744170413345e+17, 1.288744170452407e+17, 1.288744170493032e+17, 1.288744170532095e+17, 1.288744170572719e+17, 1.288744170613345e+17, 1.288744170652407e+17, 1.288744170693033e+17, 1.288744170732095e+17, 1.288744170772719e+17, 1.288744170813345e+17, 1.288744170852407e+17, 1.288744170893032e+17, 1.288744170932095e+17, 1.288744170972719e+17, 1.288744171013345e+17, 1.288744171052407e+17, 1.288744171093033e+17, 1.288744171132095e+17, 1.288744171172721e+17, 1.288744171213345e+17, 1.288744171252407e+17, 1.288744171293033e+17, 1.288744171332095e+17, 1.288744171372719e+17, 1.288744171413345e+17, 1.288744171452407e+17, 1.288744171493033e+17, 1.288744171532095e+17, 1.288744171572721e+17, 1.288744171613345e+17, 1.288744171652407e+17, 1.288744171693033e+17, 1.288744171732095e+17, 1.288744171772721e+17, 1.288744171813345e+17, 1.288744171852407e+17, 1.288744171893033e+17, 1.288744171932095e+17, 1.288744171972721e+17, 1.288744172013345e+17, 1.288744172052408e+17, 1.288744172093033e+17, 1.288744172132095e+17, 1.288744172172721e+17, 1.288744172213344e+17, 1.288744172252407e+17, 1.288744172293033e+17, 1.288744172332095e+17, 1.288744172372721e+17, 1.288744172413345e+17, 1.288744172452408e+17, 1.288744172493032e+17, 1.288744172532095e+17, 1.288744172572721e+17, 1.288744172613344e+17, 1.288744172652408e+17, 1.288744172693032e+17, 1.288744172732095e+17, 1.288744172772719e+17, 1.288744172813345e+17, 1.288744172852408e+17, 1.288744172893032e+17, 1.288744172932096e+17, 1.288744172972719e+17, 1.288744173013345e+17, 1.288744173052407e+17, 1.288744173093032e+17, 1.288744173132095e+17, 1.288744173172719e+17, 1.288744173213345e+17, 1.288744173252407e+17, 1.288744173293033e+17, 1.288744173332095e+17, 1.288744173372719e+17, 1.288744173413345e+17, 1.288744173452407e+17, 1.288744173493032e+17, 1.288744173532095e+17, 1.288744173572719e+17, 1.288744173613345e+17, 1.288744173652407e+17, 1.288744173693033e+17, 1.288744173732095e+17, 1.288744173772721e+17, 1.288744173813345e+17, 1.288744173852407e+17, 1.288744173893033e+17, 1.288744173932095e+17, 1.288744173972719e+17, 1.288744174013345e+17, 1.288744174052407e+17, 1.288744174093033e+17, 1.288744174132095e+17, 1.288744174172721e+17, 1.288744174213345e+17, 1.288744174252407e+17, 1.288744174293033e+17, 1.288744174332095e+17, 1.288744174372721e+17, 1.288744174413345e+17, 1.288744174452407e+17, 1.288744174493033e+17, 1.288744174532095e+17, 1.288744174572721e+17, 1.288744174613344e+17, 1.288744174652408e+17, 1.288744174693033e+17, 1.288744174732095e+17, 1.288744174772721e+17, 1.288744174813344e+17, 1.288744174852407e+17, 1.288744174893032e+17, 1.288744174932095e+17, 1.288744174972721e+17, 1.288744175013345e+17, 1.288744175052408e+17, 1.288744175093032e+17, 1.288744175132095e+17, 1.288744175172719e+17, 1.288744175213344e+17, 1.288744175252408e+17, 1.288744175293032e+17, 1.288744175332095e+17, 1.288744175372719e+17, 1.288744175413345e+17, 1.288744175452407e+17, 1.288744175493033e+17, 1.288744175532096e+17, 1.288744175572719e+17, 1.288744175613345e+17, 1.288744175652407e+17, 1.288744175693032e+17, 1.288744175732095e+17, 1.288744175772719e+17, 1.288744175813345e+17, 1.288744175852407e+17, 1.288744175893033e+17, 1.288744175932095e+17, 1.288744175972719e+17, 1.288744176013345e+17, 1.288744176052407e+17, 1.288744176093032e+17, 1.288744176132095e+17, 1.288744176172719e+17, 1.288744176213345e+17, 1.288744176252407e+17, 1.288744176293033e+17, 1.288744176332095e+17, 1.288744176372721e+17, 1.288744176413345e+17, 1.288744176452407e+17, 1.288744176493033e+17, 1.288744176532095e+17, 1.288744176572719e+17, 1.288744176613345e+17, 1.288744176652407e+17, 1.288744176693033e+17, 1.288744176732095e+17, 1.288744176772721e+17, 1.288744176813345e+17, 1.288744176852407e+17, 1.288744176893033e+17, 1.288744176932095e+17, 1.288744176972721e+17, 1.288744177013345e+17, 1.288744177052407e+17, 1.288744177093033e+17, 1.288744177132095e+17, 1.288744177172721e+17, 1.288744177213344e+17, 1.288744177252408e+17, 1.288744177293033e+17, 1.288744177332095e+17, 1.288744177372721e+17, 1.288744177413344e+17, 1.288744177452407e+17, 1.288744177493032e+17, 1.288744177532095e+17, 1.288744177572721e+17, 1.288744177613345e+17, 1.288744177652408e+17, 1.288744177693032e+17, 1.288744177732096e+17, 1.288744177772719e+17, 1.288744177813344e+17, 1.288744177852408e+17, 1.288744177893032e+17, 1.288744177932095e+17, 1.288744177972719e+17, 1.288744178013345e+17, 1.288744178052407e+17, 1.288744178093033e+17, 1.288744178132096e+17, 1.288744178172719e+17, 1.288744178213345e+17, 1.288744178252407e+17, 1.288744178293032e+17, 1.288744178332095e+17, 1.288744178372719e+17, 1.288744178413345e+17, 1.288744178452407e+17, 1.288744178493033e+17, 1.288744178532095e+17, 1.288744178572719e+17, 1.288744178613345e+17, 1.288744178652407e+17, 1.288744178693033e+17, 1.288744178732095e+17, 1.288744178772719e+17, 1.288744178813345e+17, 1.288744178852407e+17, 1.288744178893033e+17, 1.288744178932095e+17, 1.288744178972721e+17, 1.288744179013345e+17, 1.288744179052407e+17, 1.288744179093033e+17, 1.288744179132095e+17, 1.288744179172719e+17, 1.288744179213345e+17, 1.288744179252407e+17, 1.288744179293033e+17, 1.288744179332095e+17, 1.288744179372721e+17, 1.288744179413345e+17, 1.288744179452407e+17, 1.288744179493033e+17, 1.288744179532095e+17, 1.288744179572721e+17, 1.288744179613345e+17, 1.288744179652407e+17, 1.288744179693033e+17, 1.288744179732095e+17, 1.288744179772721e+17, 1.288744179813344e+17, 1.288744179852408e+17, 1.288744179893033e+17, 1.288744179932095e+17, 1.288744179972721e+17, 1.288744180013344e+17, 1.288744180052407e+17, 1.288744180093032e+17, 1.288744180132095e+17, 1.288744180172721e+17, 1.288744180213345e+17, 1.288744180252408e+17, 1.288744180293032e+17, 1.288744180332096e+17, 1.288744180372719e+17, 1.288744180413344e+17, 1.288744180452408e+17, 1.288744180493032e+17, 1.288744180532095e+17, 1.288744180572719e+17, 1.288744180613345e+17, 1.288744180652407e+17, 1.288744180693033e+17, 1.288744180732096e+17, 1.288744180772719e+17, 1.288744180813345e+17, 1.288744180852407e+17, 1.288744180893032e+17, 1.288744180932095e+17, 1.288744180972719e+17, 1.288744181013345e+17, 1.288744181052407e+17, 1.288744181093033e+17, 1.288744181132095e+17, 1.288744181172719e+17, 1.288744181213345e+17, 1.288744181252407e+17, 1.288744181293033e+17, 1.288744181332095e+17, 1.288744181372719e+17, 1.288744181413345e+17, 1.288744181452407e+17, 1.288744181493033e+17, 1.288744181532095e+17, 1.288744181572721e+17, 1.288744181613345e+17, 1.288744181652407e+17, 1.288744181693033e+17, 1.288744181732095e+17, 1.288744181772719e+17, 1.288744181813345e+17, 1.288744181852407e+17, 1.288744181893033e+17, 1.288744181932095e+17, 1.288744181972721e+17, 1.288744182013345e+17, 1.288744182052407e+17, 1.288744182093033e+17, 1.288744182132095e+17, 1.288744182172721e+17, 1.288744182213345e+17, 1.288744182252407e+17, 1.288744182293033e+17, 1.288744182332095e+17, 1.288744182372721e+17, 1.288744182413345e+17, 1.288744182452408e+17, 1.288744182493033e+17, 1.288744182532095e+17, 1.288744182572721e+17, 1.288744182613344e+17, 1.288744182652407e+17, 1.288744182693032e+17, 1.288744182732095e+17, 1.288744182772721e+17, 1.288744182813345e+17, 1.288744182852408e+17, 1.288744182893032e+17, 1.288744182932096e+17, 1.288744182972719e+17, 1.288744183013344e+17, 1.288744183052408e+17, 1.288744183093032e+17, 1.288744183132095e+17, 1.288744183172719e+17, 1.288744183213345e+17, 1.288744183252407e+17, 1.288744183293033e+17, 1.288744183332096e+17, 1.288744183372719e+17, 1.288744183413345e+17, 1.288744183452407e+17, 1.288744183493032e+17, 1.288744183532095e+17, 1.288744183572719e+17, 1.288744183613345e+17, 1.288744183652407e+17, 1.288744183693033e+17, 1.288744183732095e+17, 1.288744183772719e+17, 1.288744183813345e+17, 1.288744183852407e+17, 1.288744183893033e+17, 1.288744183932095e+17, 1.288744183972719e+17, 1.288744184013345e+17, 1.288744184052407e+17, 1.288744184093033e+17, 1.288744184132095e+17, 1.288744184172721e+17, 1.288744184213345e+17, 1.288744184252407e+17, 1.288744184293033e+17, 1.288744184332095e+17, 1.288744184372719e+17, 1.288744184413345e+17, 1.288744184452407e+17, 1.288744184493033e+17, 1.288744184532095e+17, 1.288744184572721e+17, 1.288744184613345e+17, 1.288744184652408e+17, 1.288744184693033e+17, 1.288744184732095e+17, 1.288744184772721e+17, 1.288744184813344e+17, 1.288744184852407e+17, 1.288744184893033e+17, 1.288744184932095e+17, 1.288744184972721e+17, 1.288744185013345e+17, 1.288744185052408e+17, 1.288744185093032e+17, 1.288744185132095e+17, 1.288744185172721e+17, 1.288744185213344e+17, 1.288744185252408e+17, 1.288744185293032e+17, 1.288744185332095e+17, 1.288744185372719e+17, 1.288744185413345e+17, 1.288744185452408e+17, 1.288744185493032e+17, 1.288744185532096e+17, 1.288744185572719e+17, 1.288744185613345e+17, 1.288744185652407e+17, 1.288744185693032e+17, 1.288744185732095e+17, 1.288744185772719e+17, 1.288744185813345e+17, 1.288744185852407e+17, 1.288744185893033e+17, 1.288744185932095e+17, 1.288744185972719e+17, 1.288744186013345e+17, 1.288744186052407e+17, 1.288744186093032e+17, 1.288744186132095e+17, 1.288744186172719e+17, 1.288744186213345e+17, 1.288744186252407e+17, 1.288744186293033e+17, 1.288744186332095e+17, 1.288744186372719e+17, 1.288744186413345e+17, 1.288744186452407e+17, 1.288744186493033e+17, 1.288744186532095e+17, 1.288744186572719e+17, 1.288744186613345e+17, 1.288744186652407e+17, 1.288744186693033e+17, 1.288744186732095e+17, 1.288744186772721e+17, 1.288744186813345e+17, 1.288744186852407e+17, 1.288744186893033e+17, 1.288744186932095e+17, 1.288744186972719e+17, 1.288744187013345e+17, 1.288744187052407e+17, 1.288744187093033e+17, 1.288744187132095e+17, 1.288744187172721e+17, 1.288744187213345e+17, 1.288744187252408e+17, 1.288744187293033e+17, 1.288744187332095e+17, 1.288744187372721e+17, 1.288744187413344e+17, 1.288744187452407e+17, 1.288744187493033e+17, 1.288744187532095e+17, 1.288744187572721e+17, 1.288744187613345e+17, 1.288744187652408e+17, 1.288744187693032e+17, 1.288744187732095e+17, 1.288744187772721e+17, 1.288744187813344e+17, 1.288744187852408e+17, 1.288744187893032e+17, 1.288744187932095e+17, 1.288744187972719e+17, 1.288744188013345e+17, 1.288744188052408e+17, 1.288744188093032e+17, 1.288744188132096e+17, 1.288744188172719e+17, 1.288744188213345e+17, 1.288744188252407e+17, 1.288744188293032e+17, 1.288744188332095e+17, 1.288744188372719e+17, 1.288744188413345e+17, 1.288744188452407e+17, 1.288744188493033e+17, 1.288744188532095e+17, 1.288744188572719e+17, 1.288744188613345e+17, 1.288744188652407e+17, 1.288744188693032e+17, 1.288744188732095e+17, 1.288744188772719e+17, 1.288744188813345e+17, 1.288744188852407e+17, 1.288744188893033e+17, 1.288744188932095e+17, 1.288744188972721e+17, 1.288744189013345e+17, 1.288744189052407e+17, 1.288744189093033e+17, 1.288744189132095e+17, 1.288744189172719e+17, 1.288744189213345e+17, 1.288744189252407e+17, 1.288744189293033e+17, 1.288744189332095e+17, 1.288744189372721e+17, 1.288744189413345e+17, 1.288744189452407e+17, 1.288744189493033e+17, 1.288744189532095e+17, 1.288744189572719e+17, 1.288744189613345e+17, 1.288744189652407e+17, 1.288744189693033e+17, 1.288744189732095e+17, 1.288744189772721e+17, 1.288744189813345e+17, 1.288744189852408e+17, 1.288744189893033e+17, 1.288744189932095e+17, 1.288744189972721e+17, 1.288744190013344e+17, 1.288744190052407e+17, 1.288744190093033e+17, 1.288744190132095e+17, 1.288744190172721e+17, 1.288744190213345e+17, 1.288744190252408e+17, 1.288744190293032e+17, 1.288744190332095e+17, 1.288744190372721e+17, 1.288744190413344e+17, 1.288744190452408e+17, 1.288744190493032e+17, 1.288744190532095e+17, 1.288744190572719e+17, 1.288744190613345e+17, 1.288744190652408e+17, 1.288744190693032e+17, 1.288744190732096e+17, 1.288744190772719e+17, 1.288744190813345e+17, 1.288744190852407e+17, 1.288744190893032e+17, 1.288744190932095e+17, 1.288744190972719e+17, 1.288744191013345e+17, 1.288744191052407e+17, 1.288744191093033e+17, 1.288744191132095e+17, 1.288744191172719e+17, 1.288744191213345e+17, 1.288744191252407e+17, 1.288744191293032e+17, 1.288744191332095e+17, 1.288744191372719e+17, 1.288744191413345e+17, 1.288744191452407e+17, 1.288744191493033e+17, 1.288744191532095e+17, 1.288744191572721e+17, 1.288744191613345e+17, 1.288744191652407e+17, 1.288744191693033e+17, 1.288744191732095e+17, 1.288744191772719e+17, 1.288744191813345e+17, 1.288744191852407e+17, 1.288744191893033e+17, 1.288744191932095e+17, 1.288744191972721e+17, 1.288744192013345e+17, 1.288744192052407e+17, 1.288744192093033e+17, 1.288744192132095e+17, 1.288744192172721e+17, 1.288744192213345e+17, 1.288744192252407e+17, 1.288744192293033e+17, 1.288744192332095e+17, 1.288744192372721e+17, 1.288744192413345e+17, 1.288744192452408e+17, 1.288744192493033e+17, 1.288744192532095e+17, 1.288744192572721e+17, 1.288744192613344e+17, 1.288744192652407e+17, 1.288744192693033e+17, 1.288744192732095e+17, 1.288744192772721e+17, 1.288744192813345e+17, 1.288744192852408e+17, 1.288744192893032e+17, 1.288744192932095e+17, 1.288744192972721e+17, 1.288744193013344e+17, 1.288744193052408e+17, 1.288744193093032e+17, 1.288744193132095e+17, 1.288744193172719e+17, 1.288744193213345e+17, 1.288744193252408e+17, 1.288744193293032e+17, 1.288744193332096e+17, 1.288744193372719e+17, 1.288744193413345e+17, 1.288744193452407e+17, 1.288744193493032e+17, 1.288744193532095e+17, 1.288744193572719e+17, 1.288744193613345e+17, 1.288744193652407e+17, 1.288744193693033e+17, 1.288744193732095e+17, 1.288744193772719e+17, 1.288744193813345e+17, 1.288744193852407e+17, 1.288744193893032e+17, 1.288744193932095e+17, 1.288744193972719e+17, 1.288744194013345e+17, 1.288744194052407e+17, 1.288744194093033e+17, 1.288744194132095e+17, 1.288744194172721e+17, 1.288744194213345e+17, 1.288744194252407e+17, 1.288744194293033e+17, 1.288744194332095e+17, 1.288744194372719e+17, 1.288744194413345e+17, 1.288744194452407e+17, 1.288744194493033e+17, 1.288744194532095e+17, 1.288744194572721e+17, 1.288744194613345e+17, 1.288744194652407e+17, 1.288744194693033e+17, 1.288744194732095e+17, 1.288744194772721e+17, 1.288744194813345e+17, 1.288744194852407e+17, 1.288744194893033e+17, 1.288744194932095e+17, 1.288744194972721e+17, 1.288744195013344e+17, 1.288744195052408e+17, 1.288744195093033e+17, 1.288744195132095e+17, 1.288744195172721e+17, 1.288744195213344e+17, 1.288744195252407e+17, 1.288744195293032e+17, 1.288744195332095e+17, 1.288744195372721e+17, 1.288744195413345e+17, 1.288744195452408e+17, 1.288744195493032e+17, 1.288744195532096e+17, 1.288744195572719e+17, 1.288744195613344e+17, 1.288744195652408e+17, 1.288744195693032e+17, 1.288744195732095e+17, 1.288744195772719e+17, 1.288744195813345e+17, 1.288744195852407e+17, 1.288744195893033e+17, 1.288744195932096e+17, 1.288744195972719e+17, 1.288744196013345e+17, 1.288744196052407e+17, 1.288744196093032e+17, 1.288744196132095e+17, 1.288744196172719e+17, 1.288744196213345e+17, 1.288744196252407e+17, 1.288744196293033e+17, 1.288744196332095e+17, 1.288744196372719e+17, 1.288744196413345e+17, 1.288744196452407e+17, 1.288744196493032e+17, 1.288744196532095e+17, 1.288744196572719e+17, 1.288744196613345e+17, 1.288744196652407e+17, 1.288744196693033e+17, 1.288744196732095e+17, 1.288744196772721e+17, 1.288744196813345e+17, 1.288744196852407e+17, 1.288744196893033e+17, 1.288744196932095e+17, 1.288744196972719e+17, 1.288744197013345e+17, 1.288744197052407e+17, 1.288744197093033e+17, 1.288744197132095e+17, 1.288744197172721e+17, 1.288744197213345e+17, 1.288744197252407e+17, 1.288744197293033e+17, 1.288744197332095e+17, 1.288744197372721e+17, 1.288744197413345e+17, 1.288744197452407e+17, 1.288744197493033e+17, 1.288744197532095e+17, 1.288744197572721e+17, 1.288744197613344e+17, 1.288744197652408e+17, 1.288744197693033e+17, 1.288744197732095e+17, 1.288744197772721e+17, 1.288744197813344e+17, 1.288744197852407e+17, 1.288744197893032e+17, 1.288744197932095e+17, 1.288744197972721e+17, 1.288744198013345e+17, 1.288744198052408e+17, 1.288744198093032e+17, 1.288744198132096e+17, 1.288744198172719e+17, 1.288744198213344e+17, 1.288744198252408e+17, 1.288744198293032e+17, 1.288744198332095e+17, 1.288744198372719e+17, 1.288744198413345e+17, 1.288744198452407e+17, 1.288744198493033e+17, 1.288744198532096e+17, 1.288744198572719e+17, 1.288744198613345e+17, 1.288744198652407e+17, 1.288744198693032e+17, 1.288744198732095e+17, 1.288744198772719e+17, 1.288744198813345e+17, 1.288744198852407e+17, 1.288744198893033e+17, 1.288744198932095e+17, 1.288744198972719e+17, 1.288744199013345e+17, 1.288744199052407e+17, 1.288744199093033e+17, 1.288744199132095e+17, 1.288744199172719e+17, 1.288744199213345e+17, 1.288744199252407e+17, 1.288744199293033e+17, 1.288744199332095e+17, 1.288744199372721e+17, 1.288744199413345e+17, 1.288744199452407e+17, 1.288744199493033e+17, 1.288744199532095e+17, 1.288744199572719e+17, 1.288744199613345e+17, 1.288744199652407e+17, 1.288744199693033e+17, 1.288744199732095e+17, 1.288744199772721e+17, 1.288744199813345e+17, 1.288744199852407e+17, 1.288744199893033e+17, 1.288744199932095e+17, 1.288744199972721e+17, 1.288744200013345e+17, 1.288744200052407e+17, 1.288744200093033e+17, 1.288744200132095e+17, 1.288744200172721e+17, 1.288744200213344e+17, 1.288744200252408e+17, 1.288744200293033e+17, 1.288744200332095e+17, 1.288744200372721e+17, 1.288744200413344e+17, 1.288744200452407e+17, 1.288744200493032e+17, 1.288744200532095e+17, 1.288744200572721e+17, 1.288744200613345e+17, 1.288744200652408e+17, 1.288744200693032e+17, 1.288744200732096e+17, 1.288744200772719e+17, 1.288744200813344e+17, 1.288744200852408e+17, 1.288744200893032e+17, 1.288744200932095e+17, 1.288744200972719e+17, 1.288744201013345e+17, 1.288744201052407e+17, 1.288744201093033e+17, 1.288744201132096e+17, 1.288744201172719e+17, 1.288744201213345e+17, 1.288744201252407e+17, 1.288744201293032e+17, 1.288744201332095e+17, 1.288744201372719e+17, 1.288744201413345e+17, 1.288744201452407e+17, 1.288744201493033e+17, 1.288744201532095e+17, 1.288744201572719e+17, 1.288744201613345e+17, 1.288744201652407e+17, 1.288744201693033e+17, 1.288744201732095e+17, 1.288744201772719e+17, 1.288744201813345e+17, 1.288744201852407e+17, 1.288744201894595e+17, 1.288744201932095e+17, 1.288744201972721e+17, 1.288744202013345e+17, 1.288744202052407e+17, 1.288744202094595e+17, 1.288744202133658e+17, 1.288744202175845e+17, 1.288744202214908e+17, 1.28874420225397e+17, 1.288744202293033e+17, 1.288744202332095e+17, 1.288744202372721e+17, 1.288744202413345e+17, 1.288744202452408e+17, 1.288744202493033e+17, 1.288744202532095e+17, 1.288744202572721e+17, 1.288744202613344e+17, 1.288744202652407e+17, 1.288744202693033e+17, 1.288744202732095e+17, 1.288744202772721e+17, 1.288744202813345e+17, 1.288744202852408e+17, 1.288744202893032e+17, 1.288744202932095e+17, 1.288744202972721e+17, 1.288744203013344e+17, 1.288744203052407e+17, 1.288744203093032e+17, 1.288744203132095e+17, 1.288744203172721e+17, 1.288744203213345e+17, 1.288744203252408e+17, 1.288744203293032e+17, 1.288744203332096e+17, 1.288744203372719e+17, 1.288744203413345e+17, 1.288744203452408e+17, 1.288744203493032e+17, 1.288744203532095e+17, 1.288744203572719e+17, 1.288744203613345e+17, 1.288744203652407e+17, 1.288744203693033e+17, 1.288744203732096e+17, 1.288744203772719e+17, 1.288744203813345e+17, 1.288744203852407e+17, 1.288744203893032e+17, 1.288744203932095e+17, 1.288744203972719e+17, 1.288744204013345e+17, 1.288744204052407e+17, 1.288744204093033e+17, 1.288744204132095e+17, 1.288744204172719e+17, 1.288744204213345e+17, 1.288744204252407e+17, 1.288744204293033e+17, 1.288744204332095e+17, 1.288744204372719e+17, 1.288744204413345e+17, 1.288744204452407e+17, 1.288744204493033e+17, 1.288744204532095e+17, 1.288744204572721e+17, 1.288744204613345e+17, 1.288744204652407e+17, 1.288744204693033e+17, 1.288744204732095e+17, 1.288744204772719e+17, 1.288744204813345e+17, 1.288744204852407e+17, 1.288744204893033e+17, 1.288744204932095e+17, 1.288744204972721e+17, 1.288744205013345e+17, 1.288744205052408e+17, 1.288744205093033e+17, 1.288744205132095e+17, 1.288744205172721e+17, 1.288744205213344e+17, 1.288744205252407e+17, 1.288744205293033e+17, 1.288744205332095e+17, 1.288744205372721e+17, 1.288744205413345e+17, 1.288744205452408e+17, 1.288744205493032e+17, 1.288744205532095e+17, 1.288744205572721e+17, 1.288744205613344e+17, 1.288744205652408e+17, 1.288744205693032e+17, 1.288744205732095e+17, 1.288744205772719e+17, 1.288744205813345e+17, 1.288744205852408e+17, 1.288744205893032e+17, 1.288744205932096e+17, 1.288744205972719e+17, 1.288744206013345e+17, 1.288744206052407e+17, 1.288744206093032e+17, 1.288744206132095e+17, 1.288744206172719e+17, 1.288744206213345e+17, 1.288744206252407e+17, 1.288744206293033e+17, 1.288744206332095e+17, 1.288744206372719e+17, 1.288744206413345e+17, 1.288744206452407e+17, 1.288744206493032e+17, 1.288744206532095e+17, 1.288744206572719e+17, 1.288744206613345e+17, 1.288744206652407e+17, 1.288744206693033e+17, 1.288744206732095e+17, 1.288744206772719e+17, 1.288744206813345e+17, 1.288744206852407e+17, 1.288744206893033e+17, 1.288744206932095e+17, 1.288744206972719e+17, 1.288744207013345e+17, 1.288744207052407e+17, 1.288744207093033e+17, 1.288744207132095e+17, 1.288744207172721e+17, 1.288744207213345e+17, 1.288744207252407e+17, 1.288744207293033e+17, 1.288744207332095e+17, 1.288744207372719e+17, 1.288744207413345e+17, 1.288744207452407e+17, 1.288744207493033e+17, 1.288744207532095e+17, 1.288744207572721e+17, 1.288744207613345e+17, 1.288744207652408e+17, 1.288744207693033e+17, 1.288744207732095e+17, 1.288744207772721e+17, 1.288744207813344e+17, 1.288744207852407e+17, 1.288744207893033e+17, 1.288744207932095e+17, 1.288744207972721e+17, 1.288744208013345e+17, 1.288744208052408e+17, 1.288744208093032e+17, 1.288744208132095e+17, 1.288744208172721e+17, 1.288744208213344e+17, 1.288744208252408e+17, 1.288744208293032e+17, 1.288744208332095e+17, 1.288744208372719e+17, 1.288744208413345e+17, 1.288744208452408e+17, 1.288744208493032e+17, 1.288744208532096e+17, 1.288744208572719e+17, 1.288744208613345e+17, 1.288744208652407e+17, 1.288744208693032e+17, 1.288744208732095e+17, 1.288744208772719e+17, 1.288744208813345e+17, 1.288744208852407e+17, 1.288744208893033e+17, 1.288744208932095e+17, 1.288744208972719e+17, 1.288744209013345e+17, 1.288744209052407e+17, 1.288744209093032e+17, 1.288744209132095e+17, 1.288744209172719e+17, 1.288744209213345e+17, 1.288744209252407e+17, 1.288744209293033e+17, 1.288744209332095e+17, 1.288744209372721e+17, 1.288744209413345e+17, 1.288744209452407e+17, 1.288744209493033e+17, 1.288744209532095e+17, 1.288744209572719e+17, 1.288744209613345e+17, 1.288744209652407e+17, 1.288744209693033e+17, 1.288744209732095e+17, 1.288744209772721e+17, 1.288744209813345e+17, 1.288744209852407e+17, 1.288744209893033e+17, 1.288744209932095e+17, 1.288744209972721e+17, 1.288744210013345e+17, 1.288744210052407e+17, 1.288744210093033e+17, 1.288744210132095e+17, 1.288744210172721e+17, 1.288744210213345e+17, 1.288744210252408e+17, 1.288744210293033e+17, 1.288744210332095e+17, 1.288744210372721e+17, 1.288744210413344e+17, 1.288744210452407e+17, 1.288744210493033e+17, 1.288744210532095e+17, 1.288744210572721e+17, 1.288744210613345e+17, 1.288744210652408e+17, 1.288744210693032e+17, 1.288744210732095e+17, 1.288744210772721e+17, 1.288744210813344e+17, 1.288744210852408e+17, 1.288744210893032e+17, 1.288744210932095e+17, 1.288744210972719e+17, 1.288744211013345e+17, 1.288744211052408e+17, 1.288744211093032e+17, 1.288744211132096e+17, 1.288744211172719e+17, 1.288744211213345e+17, 1.288744211252407e+17, 1.288744211293032e+17, 1.288744211332095e+17, 1.288744211372719e+17, 1.288744211413345e+17, 1.288744211452407e+17, 1.288744211493033e+17, 1.288744211532095e+17, 1.288744211572719e+17, 1.288744211613345e+17, 1.288744211652407e+17, 1.288744211693032e+17, 1.288744211732095e+17, 1.288744211772719e+17, 1.288744211813345e+17, 1.288744211852407e+17, 1.288744211893033e+17, 1.288744211932095e+17, 1.288744211972721e+17, 1.288744212013345e+17, 1.288744212052407e+17, 1.288744212093033e+17, 1.288744212132095e+17, 1.288744212172719e+17, 1.288744212213345e+17, 1.288744212252407e+17, 1.288744212293033e+17, 1.288744212332095e+17, 1.288744212372721e+17, 1.288744212413345e+17, 1.288744212452407e+17, 1.288744212493033e+17, 1.288744212532095e+17, 1.288744212572721e+17, 1.288744212613345e+17, 1.288744212652407e+17, 1.288744212693033e+17, 1.288744212732095e+17, 1.288744212772721e+17, 1.288744212813344e+17, 1.288744212852408e+17, 1.288744212893033e+17, 1.288744212932095e+17, 1.288744212972721e+17, 1.288744213013344e+17, 1.288744213052407e+17, 1.288744213093032e+17, 1.288744213132095e+17, 1.288744213172721e+17, 1.288744213213345e+17, 1.288744213252408e+17, 1.288744213293032e+17, 1.288744213332095e+17, 1.288744213372719e+17, 1.288744213413344e+17, 1.288744213452408e+17, 1.288744213493032e+17, 1.288744213532095e+17, 1.288744213572719e+17, 1.288744213613345e+17, 1.288744213652407e+17, 1.288744213693032e+17, 1.288744213732096e+17, 1.288744213772719e+17, 1.288744213813345e+17, 1.288744213852407e+17, 1.288744213893032e+17, 1.288744213932095e+17, 1.288744213972719e+17, 1.288744214013345e+17, 1.288744214052407e+17, 1.288744214093033e+17, 1.288744214132095e+17, 1.288744214172719e+17, 1.288744214213345e+17, 1.288744214252407e+17, 1.288744214293032e+17, 1.288744214332095e+17, 1.288744214372719e+17, 1.288744214413345e+17, 1.288744214452407e+17, 1.288744214493033e+17, 1.288744214532095e+17, 1.288744214572721e+17, 1.288744214613345e+17, 1.288744214652407e+17, 1.288744214693033e+17, 1.288744214732095e+17, 1.288744214772719e+17, 1.288744214813345e+17, 1.288744214852407e+17, 1.288744214893033e+17, 1.288744214932095e+17, 1.288744214972721e+17, 1.288744215013345e+17, 1.288744215052407e+17, 1.288744215093033e+17, 1.288744215132095e+17, 1.288744215172721e+17, 1.288744215213345e+17, 1.288744215252407e+17, 1.288744215293033e+17, 1.288744215332095e+17, 1.288744215372721e+17, 1.288744215413344e+17, 1.288744215452408e+17, 1.288744215493033e+17, 1.288744215532095e+17, 1.288744215572721e+17, 1.288744215613344e+17, 1.288744215652407e+17, 1.288744215693032e+17, 1.288744215732095e+17, 1.288744215772721e+17, 1.288744215813345e+17, 1.288744215852408e+17, 1.288744215893032e+17, 1.288744215932096e+17, 1.288744215972719e+17, 1.288744216013344e+17, 1.288744216052408e+17, 1.288744216093032e+17, 1.288744216132095e+17, 1.288744216172719e+17, 1.288744216213345e+17, 1.288744216252407e+17, 1.288744216293033e+17, 1.288744216332096e+17, 1.288744216372719e+17, 1.288744216413345e+17, 1.288744216452407e+17, 1.288744216493032e+17, 1.288744216532095e+17, 1.288744216572719e+17, 1.288744216613345e+17, 1.288744216652407e+17, 1.288744216693033e+17, 1.288744216732095e+17, 1.288744216772719e+17, 1.288744216813345e+17, 1.288744216852407e+17, 1.288744216893033e+17, 1.288744216932095e+17, 1.288744216972719e+17, 1.288744217013345e+17, 1.288744217052407e+17, 1.288744217093033e+17, 1.288744217132095e+17, 1.288744217172721e+17, 1.288744217213345e+17, 1.288744217252407e+17, 1.288744217293033e+17, 1.288744217332095e+17, 1.288744217372719e+17, 1.288744217413345e+17, 1.288744217452407e+17, 1.288744217493033e+17, 1.288744217532095e+17, 1.288744217572721e+17, 1.288744217613345e+17, 1.288744217652407e+17, 1.288744217693033e+17, 1.288744217732095e+17, 1.288744217772721e+17, 1.288744217813345e+17, 1.288744217852407e+17, 1.288744217893033e+17, 1.288744217932095e+17, 1.288744217972721e+17, 1.288744218013344e+17, 1.288744218052408e+17, 1.288744218093033e+17, 1.288744218132095e+17, 1.288744218172721e+17, 1.288744218213344e+17, 1.288744218252407e+17, 1.288744218293032e+17, 1.288744218332095e+17, 1.288744218372721e+17, 1.288744218413345e+17, 1.288744218452408e+17, 1.288744218493032e+17, 1.288744218532096e+17, 1.288744218572719e+17, 1.288744218613344e+17, 1.288744218652408e+17, 1.288744218693032e+17, 1.288744218732095e+17, 1.288744218772719e+17, 1.288744218813345e+17, 1.288744218852407e+17, 1.288744218893033e+17, 1.288744218932096e+17, 1.288744218972719e+17, 1.288744219013345e+17, 1.288744219052407e+17, 1.288744219093032e+17, 1.288744219132095e+17, 1.288744219172719e+17, 1.288744219213345e+17, 1.288744219252407e+17, 1.288744219293033e+17, 1.288744219332095e+17, 1.288744219372719e+17, 1.288744219413345e+17, 1.288744219452407e+17, 1.288744219493033e+17, 1.288744219532095e+17, 1.288744219572719e+17, 1.288744219613345e+17, 1.288744219652407e+17, 1.288744219693033e+17, 1.288744219732095e+17, 1.288744219772721e+17, 1.288744219813345e+17, 1.288744219852407e+17, 1.288744219893033e+17, 1.288744219932095e+17, 1.288744219972719e+17, 1.288744220013345e+17, 1.288744220052407e+17, 1.288744220093033e+17, 1.288744220132095e+17, 1.288744220172721e+17, 1.288744220213345e+17, 1.288744220252407e+17, 1.288744220293033e+17, 1.288744220332095e+17, 1.288744220372721e+17, 1.288744220413345e+17, 1.288744220452407e+17, 1.288744220493033e+17, 1.288744220532095e+17, 1.288744220572721e+17, 1.288744220613345e+17, 1.288744220652408e+17, 1.288744220693033e+17, 1.288744220732095e+17, 1.288744220772721e+17, 1.288744220813344e+17, 1.288744220852407e+17, 1.288744220893032e+17, 1.288744220932095e+17, 1.288744220972721e+17, 1.288744221013345e+17, 1.288744221052408e+17, 1.288744221093032e+17, 1.288744221132096e+17, 1.288744221172719e+17, 1.288744221213344e+17, 1.288744221252408e+17, 1.288744221293032e+17, 1.288744221332095e+17, 1.288744221372719e+17, 1.288744221413345e+17, 1.288744221452407e+17, 1.288744221493033e+17, 1.288744221532096e+17, 1.288744221572719e+17, 1.288744221613345e+17, 1.288744221652407e+17, 1.288744221693032e+17, 1.288744221732095e+17, 1.288744221772719e+17, 1.288744221813345e+17, 1.288744221852407e+17, 1.288744221893033e+17, 1.288744221932095e+17, 1.288744221972719e+17, 1.288744222013345e+17, 1.288744222052407e+17, 1.288744222093033e+17, 1.288744222132095e+17, 1.288744222172719e+17, 1.288744222213345e+17, 1.288744222252407e+17, 1.288744222293033e+17, 1.288744222332095e+17, 1.288744222372721e+17, 1.288744222413345e+17, 1.288744222452407e+17, 1.288744222493033e+17, 1.288744222532095e+17, 1.288744222572719e+17, 1.288744222613345e+17, 1.288744222652407e+17, 1.288744222693033e+17, 1.288744222732095e+17, 1.288744222772721e+17, 1.288744222813345e+17, 1.288744222852408e+17, 1.288744222893033e+17, 1.288744222932095e+17, 1.288744222972721e+17, 1.288744223013344e+17, 1.288744223052407e+17, 1.288744223093033e+17, 1.288744223132095e+17, 1.288744223172721e+17, 1.288744223213345e+17, 1.288744223252408e+17, 1.288744223293032e+17, 1.288744223332095e+17, 1.288744223372721e+17, 1.288744223413344e+17, 1.288744223452408e+17, 1.288744223493032e+17, 1.288744223532095e+17, 1.288744223572719e+17, 1.288744223613345e+17, 1.288744223652408e+17, 1.288744223693032e+17, 1.288744223732096e+17, 1.288744223772719e+17, 1.288744223813345e+17, 1.288744223852407e+17, 1.288744223893032e+17, 1.288744223932095e+17, 1.288744223972719e+17, 1.288744224013345e+17, 1.288744224052407e+17, 1.288744224093033e+17, 1.288744224132095e+17, 1.288744224172719e+17, 1.288744224213345e+17, 1.288744224252407e+17, 1.288744224293032e+17, 1.288744224332095e+17, 1.288744224372719e+17, 1.288744224413345e+17, 1.288744224452407e+17, 1.288744224493033e+17, 1.288744224532095e+17, 1.288744224572719e+17, 1.288744224613345e+17, 1.288744224652407e+17, 1.288744224693033e+17, 1.288744224732095e+17, 1.288744224772719e+17, 1.288744224813345e+17, 1.288744224852407e+17, 1.288744224893033e+17, 1.288744224932095e+17, 1.288744224972721e+17, 1.288744225013345e+17, 1.288744225052407e+17, 1.288744225093033e+17, 1.288744225132095e+17, 1.288744225172719e+17, 1.288744225213345e+17, 1.288744225252407e+17, 1.288744225293033e+17, 1.288744225332095e+17, 1.288744225372721e+17, 1.288744225413345e+17, 1.288744225452408e+17, 1.288744225493033e+17, 1.288744225532095e+17, 1.288744225572721e+17, 1.288744225613344e+17, 1.288744225652407e+17, 1.288744225693033e+17, 1.288744225732095e+17, 1.288744225772721e+17, 1.288744225813345e+17, 1.288744225852408e+17, 1.288744225893032e+17, 1.288744225932095e+17, 1.288744225972721e+17, 1.288744226013344e+17, 1.288744226052408e+17, 1.288744226093032e+17, 1.288744226132095e+17, 1.288744226172719e+17, 1.288744226213345e+17, 1.288744226252408e+17, 1.288744226293032e+17, 1.288744226332096e+17, 1.288744226372719e+17, 1.288744226413345e+17, 1.288744226452407e+17, 1.288744226493032e+17, 1.288744226532095e+17, 1.288744226572719e+17, 1.288744226613345e+17, 1.288744226652407e+17, 1.288744226693033e+17, 1.288744226732095e+17, 1.288744226772719e+17, 1.288744226813345e+17, 1.288744226852407e+17, 1.288744226893032e+17, 1.288744226932095e+17, 1.288744226972719e+17, 1.288744227013345e+17, 1.288744227052407e+17, 1.288744227093033e+17, 1.288744227132095e+17, 1.288744227172721e+17, 1.288744227213345e+17, 1.288744227252407e+17, 1.288744227293033e+17, 1.288744227332095e+17, 1.288744227372719e+17, 1.288744227413345e+17, 1.288744227452407e+17, 1.288744227493033e+17, 1.288744227532095e+17, 1.288744227572721e+17, 1.288744227613345e+17, 1.288744227652407e+17, 1.288744227693033e+17, 1.288744227732095e+17, 1.288744227772719e+17, 1.288744227813345e+17, 1.288744227852407e+17, 1.288744227893033e+17, 1.288744227932095e+17, 1.288744227972721e+17, 1.288744228013345e+17, 1.288744228052408e+17, 1.288744228093033e+17, 1.288744228132095e+17, 1.288744228172721e+17, 1.288744228213344e+17, 1.288744228252407e+17, 1.288744228293033e+17, 1.288744228332095e+17, 1.288744228372721e+17, 1.288744228413345e+17, 1.288744228452408e+17, 1.288744228493032e+17, 1.288744228532095e+17, 1.288744228572721e+17, 1.288744228613344e+17, 1.288744228652408e+17, 1.288744228693032e+17, 1.288744228732095e+17, 1.288744228772719e+17, 1.288744228813345e+17, 1.288744228852408e+17, 1.288744228893032e+17, 1.288744228932096e+17, 1.288744228972719e+17, 1.288744229013345e+17, 1.288744229052407e+17, 1.288744229093032e+17, 1.288744229132095e+17, 1.288744229172719e+17, 1.288744229213345e+17, 1.288744229252407e+17, 1.288744229293033e+17, 1.288744229332095e+17, 1.288744229372719e+17, 1.288744229413345e+17, 1.288744229452407e+17, 1.288744229493032e+17, 1.288744229532095e+17, 1.288744229572719e+17, 1.288744229613345e+17, 1.288744229652407e+17, 1.288744229693033e+17, 1.288744229732095e+17, 1.288744229772721e+17, 1.288744229813345e+17, 1.288744229852407e+17, 1.288744229893033e+17, 1.288744229932095e+17, 1.288744229972719e+17, 1.288744230013345e+17, 1.288744230052407e+17, 1.288744230093033e+17, 1.288744230132095e+17, 1.288744230172721e+17, 1.288744230213345e+17, 1.288744230252407e+17, 1.288744230293033e+17, 1.288744230332095e+17, 1.288744230372721e+17, 1.288744230413345e+17, 1.288744230452407e+17, 1.288744230493033e+17, 1.288744230532095e+17, 1.288744230572721e+17, 1.288744230613345e+17, 1.288744230652408e+17, 1.288744230693033e+17, 1.288744230732095e+17, 1.288744230772721e+17, 1.288744230813344e+17, 1.288744230852407e+17, 1.288744230893033e+17, 1.288744230932095e+17, 1.288744230972721e+17, 1.288744231013345e+17, 1.288744231052408e+17, 1.288744231093032e+17, 1.288744231132095e+17, 1.288744231172721e+17, 1.288744231213344e+17, 1.288744231252408e+17, 1.288744231293032e+17, 1.288744231332095e+17, 1.288744231372719e+17, 1.288744231413345e+17, 1.288744231452408e+17, 1.288744231493032e+17, 1.288744231532096e+17, 1.288744231572719e+17, 1.288744231613345e+17, 1.288744231652407e+17, 1.288744231693032e+17, 1.288744231732095e+17, 1.288744231772719e+17, 1.288744231813345e+17, 1.288744231852407e+17, 1.288744231893033e+17, 1.288744231932095e+17, 1.288744231972719e+17, 1.288744232013345e+17, 1.288744232052407e+17, 1.288744232093032e+17, 1.288744232132095e+17, 1.288744232172719e+17, 1.288744232213345e+17, 1.288744232252407e+17, 1.288744232293033e+17, 1.288744232332095e+17, 1.288744232372721e+17, 1.288744232413345e+17, 1.288744232452407e+17, 1.288744232493033e+17, 1.288744232532095e+17, 1.288744232572719e+17, 1.288744232613345e+17, 1.288744232652407e+17, 1.288744232693033e+17, 1.288744232732095e+17, 1.288744232772721e+17, 1.288744232813345e+17, 1.288744232852407e+17, 1.288744232893033e+17, 1.288744232932095e+17, 1.288744232972721e+17, 1.288744233013345e+17, 1.288744233052407e+17, 1.288744233093033e+17, 1.288744233132095e+17, 1.288744233172721e+17, 1.288744233213344e+17, 1.288744233252408e+17, 1.288744233293033e+17, 1.288744233332095e+17, 1.288744233372721e+17, 1.288744233413344e+17, 1.288744233452407e+17, 1.288744233493032e+17, 1.288744233532095e+17, 1.288744233572721e+17, 1.288744233613345e+17, 1.288744233652408e+17, 1.288744233693032e+17, 1.288744233732095e+17, 1.288744233772719e+17, 1.288744233813344e+17, 1.288744233852408e+17, 1.288744233893032e+17, 1.288744233932095e+17, 1.288744233972719e+17, 1.288744234013345e+17, 1.288744234052407e+17, 1.288744234093033e+17, 1.288744234132096e+17, 1.288744234172719e+17, 1.288744234213345e+17, 1.288744234252407e+17, 1.288744234293032e+17, 1.288744234332095e+17, 1.288744234372719e+17, 1.288744234413345e+17, 1.288744234452407e+17, 1.288744234493033e+17, 1.288744234532095e+17, 1.288744234572719e+17, 1.288744234613345e+17, 1.288744234652407e+17, 1.288744234693032e+17, 1.288744234732095e+17, 1.288744234772719e+17, 1.288744234813345e+17, 1.288744234852407e+17, 1.288744234893033e+17, 1.288744234932095e+17, 1.288744234972721e+17, 1.288744235013345e+17, 1.288744235052407e+17, 1.288744235093033e+17, 1.288744235132095e+17, 1.288744235172719e+17, 1.288744235213345e+17, 1.288744235252407e+17, 1.288744235293033e+17, 1.288744235332095e+17, 1.288744235372721e+17, 1.288744235413345e+17, 1.288744235452407e+17, 1.288744235493033e+17, 1.288744235532095e+17, 1.288744235572721e+17, 1.288744235613345e+17, 1.288744235652407e+17, 1.288744235693033e+17, 1.288744235732095e+17, 1.288744235772721e+17, 1.288744235813344e+17, 1.288744235852408e+17, 1.288744235893033e+17, 1.288744235932095e+17, 1.288744235972721e+17, 1.288744236013344e+17, 1.288744236052407e+17, 1.288744236093032e+17, 1.288744236132095e+17, 1.288744236172721e+17, 1.288744236213345e+17, 1.288744236252408e+17, 1.288744236293032e+17, 1.288744236332096e+17, 1.288744236372719e+17, 1.288744236413344e+17, 1.288744236452408e+17, 1.288744236493032e+17, 1.288744236532095e+17, 1.288744236572719e+17, 1.288744236613345e+17, 1.288744236652407e+17, 1.288744236693033e+17, 1.288744236732096e+17, 1.288744236772719e+17, 1.288744236813345e+17, 1.288744236852407e+17, 1.288744236893032e+17, 1.288744236932095e+17, 1.288744236972719e+17, 1.288744237013345e+17, 1.288744237052407e+17, 1.288744237093033e+17, 1.288744237132095e+17, 1.288744237172719e+17, 1.288744237213345e+17, 1.288744237252407e+17, 1.288744237293033e+17, 1.288744237332095e+17, 1.288744237372719e+17, 1.288744237413345e+17, 1.288744237452407e+17, 1.288744237493033e+17, 1.288744237532095e+17, 1.288744237572721e+17, 1.288744237613345e+17, 1.288744237652407e+17, 1.288744237693033e+17, 1.288744237732095e+17, 1.288744237772719e+17, 1.288744237813345e+17, 1.288744237852407e+17, 1.288744237893033e+17, 1.288744237932095e+17, 1.288744237972721e+17, 1.288744238013345e+17, 1.288744238052407e+17, 1.288744238093033e+17, 1.288744238132095e+17, 1.288744238172721e+17, 1.288744238213345e+17, 1.288744238252407e+17, 1.288744238293033e+17, 1.288744238332095e+17, 1.288744238372721e+17, 1.288744238413344e+17, 1.288744238452408e+17, 1.288744238493033e+17, 1.288744238532095e+17, 1.288744238572721e+17, 1.288744238613344e+17, 1.288744238652407e+17, 1.288744238693032e+17, 1.288744238732095e+17, 1.288744238772721e+17, 1.288744238813345e+17, 1.288744238852408e+17, 1.288744238893032e+17, 1.288744238932096e+17, 1.288744238972719e+17, 1.288744239013344e+17, 1.288744239052408e+17, 1.288744239093032e+17, 1.288744239132095e+17, 1.288744239172719e+17, 1.288744239213345e+17, 1.288744239252407e+17, 1.288744239293033e+17, 1.288744239332096e+17, 1.288744239372719e+17, 1.288744239413345e+17, 1.288744239452407e+17, 1.288744239493032e+17, 1.288744239532095e+17, 1.288744239572719e+17, 1.288744239613345e+17, 1.288744239652407e+17, 1.288744239693033e+17, 1.288744239732095e+17, 1.288744239772719e+17, 1.288744239813345e+17, 1.288744239852407e+17, 1.288744239893033e+17, 1.288744239932095e+17, 1.288744239972719e+17, 1.288744240013345e+17, 1.288744240052407e+17, 1.288744240093033e+17, 1.288744240132095e+17, 1.288744240172721e+17, 1.288744240213345e+17, 1.288744240252407e+17, 1.288744240293033e+17, 1.288744240332095e+17, 1.288744240372719e+17, 1.288744240413345e+17, 1.288744240452407e+17, 1.288744240493033e+17, 1.288744240532095e+17, 1.288744240572721e+17, 1.288744240613345e+17, 1.288744240652408e+17, 1.288744240693033e+17, 1.288744240732095e+17, 1.288744240772721e+17, 1.288744240813345e+17, 1.288744240852407e+17, 1.288744240893033e+17, 1.288744240932095e+17, 1.288744240972721e+17, 1.288744241013345e+17, 1.288744241052408e+17, 1.288744241093033e+17, 1.288744241132095e+17, 1.288744241172721e+17, 1.288744241213344e+17, 1.288744241252407e+17, 1.288744241293032e+17, 1.288744241332095e+17, 1.288744241372721e+17, 1.288744241413345e+17, 1.288744241452408e+17, 1.288744241493032e+17, 1.288744241532096e+17, 1.288744241572719e+17, 1.288744241613345e+17, 1.288744241652408e+17, 1.288744241693032e+17, 1.288744241732095e+17, 1.288744241772719e+17, 1.288744241813345e+17, 1.288744241852407e+17, 1.288744241893033e+17, 1.288744241932096e+17, 1.288744241972719e+17, 1.288744242013345e+17, 1.288744242052407e+17, 1.288744242093032e+17, 1.288744242132095e+17, 1.288744242172719e+17, 1.288744242213345e+17, 1.288744242252407e+17, 1.288744242293033e+17, 1.288744242332095e+17, 1.288744242372719e+17, 1.288744242413345e+17, 1.288744242452407e+17, 1.288744242493033e+17, 1.288744242532095e+17, 1.288744242572719e+17, 1.288744242613345e+17, 1.288744242652407e+17, 1.288744242693033e+17, 1.288744242732095e+17, 1.288744242772721e+17, 1.288744242813345e+17, 1.288744242852407e+17, 1.288744242893033e+17, 1.288744242932095e+17, 1.288744242972719e+17, 1.288744243013345e+17, 1.288744243052407e+17, 1.288744243093033e+17, 1.288744243132095e+17, 1.288744243172721e+17, 1.288744243213345e+17, 1.288744243252408e+17, 1.288744243293033e+17, 1.288744243332095e+17, 1.288744243372721e+17, 1.288744243413344e+17, 1.288744243452407e+17, 1.288744243493033e+17, 1.288744243532095e+17, 1.288744243572721e+17, 1.288744243613345e+17, 1.288744243652408e+17, 1.288744243693032e+17, 1.288744243732095e+17, 1.288744243772721e+17, 1.288744243813344e+17, 1.288744243852408e+17, 1.288744243893032e+17, 1.288744243932095e+17, 1.288744243972719e+17, 1.288744244013345e+17, 1.288744244052408e+17, 1.288744244093032e+17, 1.288744244132096e+17, 1.288744244172719e+17, 1.288744244213345e+17, 1.288744244252407e+17, 1.288744244293032e+17, 1.288744244332095e+17, 1.288744244372719e+17, 1.288744244413345e+17, 1.288744244452407e+17, 1.288744244493033e+17, 1.288744244532095e+17, 1.288744244572719e+17, 1.288744244613345e+17, 1.288744244652407e+17, 1.288744244693032e+17, 1.288744244732095e+17, 1.288744244772719e+17, 1.288744244813345e+17, 1.288744244852407e+17, 1.288744244893033e+17, 1.288744244932095e+17, 1.288744244972719e+17, 1.288744245013345e+17, 1.288744245052407e+17, 1.288744245093033e+17, 1.288744245132095e+17, 1.288744245172719e+17, 1.288744245213345e+17, 1.288744245252407e+17, 1.288744245293033e+17, 1.288744245332095e+17, 1.288744245372721e+17, 1.288744245413345e+17, 1.288744245452407e+17, 1.288744245493033e+17, 1.288744245532095e+17, 1.288744245572719e+17, 1.288744245613345e+17, 1.288744245652407e+17, 1.288744245693033e+17, 1.288744245732095e+17, 1.288744245772721e+17, 1.288744245813345e+17, 1.288744245852408e+17, 1.288744245893033e+17, 1.288744245932095e+17, 1.288744245972721e+17, 1.288744246013344e+17, 1.288744246052407e+17, 1.288744246093033e+17, 1.288744246132095e+17, 1.288744246172721e+17, 1.288744246213345e+17, 1.288744246252408e+17, 1.288744246293032e+17, 1.288744246332095e+17, 1.288744246372721e+17, 1.288744246413344e+17, 1.288744246452408e+17, 1.288744246493032e+17, 1.288744246532095e+17, 1.288744246572719e+17, 1.288744246613345e+17, 1.288744246652408e+17, 1.288744246693032e+17, 1.288744246732096e+17, 1.288744246772719e+17, 1.288744246813345e+17, 1.288744246852407e+17, 1.288744246893032e+17, 1.288744246932095e+17, 1.288744246972719e+17, 1.288744247013345e+17, 1.288744247052407e+17, 1.288744247093033e+17, 1.288744247132095e+17, 1.288744247172719e+17, 1.288744247213345e+17, 1.288744247252407e+17, 1.288744247293032e+17, 1.288744247332095e+17, 1.288744247372719e+17, 1.288744247413345e+17, 1.288744247452407e+17, 1.288744247493033e+17, 1.288744247532095e+17, 1.288744247572721e+17, 1.288744247613345e+17, 1.288744247652407e+17, 1.288744247693033e+17, 1.288744247732095e+17, 1.288744247772719e+17, 1.288744247813345e+17, 1.288744247852407e+17, 1.288744247893033e+17, 1.288744247932095e+17, 1.288744247972721e+17, 1.288744248013345e+17, 1.288744248052407e+17, 1.288744248093033e+17, 1.288744248132095e+17, 1.288744248172719e+17, 1.288744248213345e+17, 1.288744248252407e+17, 1.288744248293033e+17, 1.288744248332095e+17, 1.288744248372721e+17, 1.288744248413345e+17, 1.288744248452408e+17, 1.288744248493033e+17, 1.288744248532095e+17, 1.288744248572721e+17, 1.288744248613344e+17, 1.288744248652407e+17, 1.288744248693033e+17, 1.288744248732095e+17, 1.288744248772721e+17, 1.288744248813345e+17, 1.288744248852408e+17, 1.288744248893032e+17, 1.288744248932095e+17, 1.288744248972721e+17, 1.288744249013344e+17, 1.288744249052408e+17, 1.288744249093032e+17, 1.288744249132095e+17, 1.288744249172719e+17, 1.288744249213345e+17, 1.288744249252408e+17, 1.288744249293032e+17, 1.288744249332096e+17, 1.288744249372719e+17, 1.288744249413345e+17, 1.288744249452407e+17, 1.288744249493032e+17, 1.288744249532095e+17, 1.288744249572719e+17, 1.288744249613345e+17, 1.288744249652407e+17, 1.288744249693033e+17, 1.288744249732095e+17, 1.288744249772719e+17, 1.288744249813345e+17, 1.288744249852407e+17, 1.288744249893032e+17, 1.288744249932095e+17, 1.288744249972719e+17, 1.288744250013345e+17, 1.288744250052407e+17, 1.288744250093033e+17, 1.288744250132095e+17, 1.288744250172721e+17, 1.288744250213345e+17, 1.288744250252407e+17, 1.288744250293033e+17, 1.288744250332095e+17, 1.288744250372719e+17, 1.288744250413345e+17, 1.288744250452407e+17, 1.288744250493033e+17, 1.288744250532095e+17, 1.288744250572721e+17, 1.288744250613345e+17, 1.288744250652407e+17, 1.288744250693033e+17, 1.288744250732095e+17, 1.288744250772721e+17, 1.288744250813345e+17, 1.288744250852407e+17, 1.288744250893033e+17, 1.288744250932095e+17, 1.288744250972721e+17, 1.288744251013344e+17, 1.288744251052408e+17, 1.288744251093033e+17, 1.288744251132095e+17, 1.288744251172721e+17, 1.288744251213344e+17, 1.288744251252407e+17, 1.288744251293032e+17, 1.288744251332095e+17, 1.288744251372721e+17, 1.288744251413345e+17, 1.288744251452408e+17, 1.288744251493032e+17, 1.288744251532095e+17, 1.288744251572719e+17, 1.288744251613344e+17, 1.288744251652408e+17, 1.288744251693032e+17, 1.288744251732095e+17, 1.288744251772719e+17, 1.288744251813345e+17, 1.288744251852407e+17, 1.288744251893032e+17, 1.288744251932096e+17, 1.288744251972719e+17, 1.288744252013345e+17, 1.288744252052407e+17, 1.288744252093032e+17, 1.288744252132095e+17, 1.288744252172719e+17, 1.288744252213345e+17, 1.288744252252407e+17, 1.288744252293033e+17, 1.288744252332095e+17, 1.288744252372719e+17, 1.288744252413345e+17, 1.288744252452407e+17, 1.288744252493032e+17, 1.288744252532095e+17, 1.288744252572719e+17, 1.288744252613345e+17, 1.288744252652407e+17, 1.288744252693033e+17, 1.288744252732095e+17, 1.288744252772721e+17, 1.288744252813345e+17, 1.288744252852407e+17, 1.288744252893033e+17, 1.288744252932095e+17, 1.288744252972719e+17, 1.288744253013345e+17, 1.288744253052407e+17, 1.288744253093033e+17, 1.288744253132095e+17, 1.288744253172721e+17, 1.288744253213345e+17, 1.288744253252407e+17, 1.288744253293033e+17, 1.288744253332095e+17, 1.288744253372721e+17, 1.288744253413345e+17, 1.288744253452407e+17, 1.288744253493033e+17, 1.288744253532095e+17, 1.288744253572721e+17, 1.288744253613344e+17, 1.288744253652408e+17, 1.288744253693033e+17, 1.288744253732095e+17, 1.288744253772721e+17, 1.288744253813344e+17, 1.288744253852407e+17, 1.288744253893032e+17, 1.288744253932095e+17, 1.288744253972721e+17, 1.288744254013345e+17, 1.288744254052408e+17, 1.288744254093032e+17, 1.288744254132096e+17, 1.288744254172719e+17, 1.288744254213344e+17, 1.288744254252408e+17, 1.288744254293032e+17, 1.288744254332095e+17, 1.288744254372719e+17, 1.288744254413345e+17, 1.288744254452407e+17, 1.288744254493033e+17, 1.288744254532096e+17, 1.288744254572719e+17, 1.288744254613345e+17, 1.288744254652407e+17, 1.288744254693032e+17, 1.288744254732095e+17, 1.288744254772719e+17, 1.288744254813345e+17, 1.288744254852407e+17, 1.288744254893033e+17, 1.288744254932095e+17, 1.288744254972719e+17, 1.288744255013345e+17, 1.288744255052407e+17, 1.288744255093033e+17, 1.288744255132095e+17, 1.288744255172719e+17, 1.288744255213345e+17, 1.288744255252407e+17, 1.288744255293033e+17, 1.288744255332095e+17, 1.288744255372721e+17, 1.288744255413345e+17, 1.288744255452407e+17, 1.288744255493033e+17, 1.288744255532095e+17, 1.288744255572719e+17, 1.288744255613345e+17, 1.288744255652407e+17, 1.288744255693033e+17, 1.288744255732095e+17, 1.288744255772721e+17, 1.288744255813345e+17, 1.288744255852407e+17, 1.288744255893033e+17, 1.288744255932095e+17, 1.288744255972721e+17, 1.288744256013345e+17, 1.288744256052407e+17, 1.288744256093033e+17, 1.288744256132095e+17, 1.288744256172721e+17, 1.288744256213344e+17, 1.288744256252408e+17, 1.288744256293033e+17, 1.288744256332095e+17, 1.288744256372721e+17, 1.288744256413344e+17, 1.288744256452407e+17, 1.288744256493032e+17, 1.288744256532095e+17, 1.288744256572721e+17, 1.288744256613345e+17, 1.288744256652408e+17, 1.288744256693032e+17, 1.288744256732096e+17, 1.288744256772719e+17, 1.288744256813344e+17, 1.288744256852408e+17, 1.288744256893032e+17, 1.288744256932095e+17, 1.288744256972719e+17, 1.288744257013345e+17, 1.288744257052407e+17, 1.288744257093033e+17, 1.288744257132096e+17, 1.288744257172719e+17, 1.288744257213345e+17, 1.288744257252407e+17, 1.288744257293032e+17, 1.288744257332095e+17, 1.288744257372719e+17, 1.288744257413345e+17, 1.288744257452407e+17, 1.288744257493033e+17, 1.288744257532095e+17, 1.288744257572719e+17, 1.288744257613345e+17, 1.288744257652407e+17, 1.288744257693033e+17, 1.288744257732095e+17, 1.288744257772719e+17, 1.288744257813345e+17, 1.288744257852407e+17, 1.288744257893033e+17, 1.288744257932095e+17, 1.288744257972721e+17, 1.288744258013345e+17, 1.288744258052407e+17, 1.288744258093033e+17, 1.288744258132095e+17, 1.288744258172719e+17, 1.288744258213345e+17, 1.288744258252407e+17, 1.288744258293033e+17, 1.288744258332095e+17, 1.288744258372721e+17, 1.288744258413345e+17, 1.288744258452407e+17, 1.288744258493033e+17, 1.288744258532095e+17, 1.288744258572721e+17, 1.288744258613345e+17, 1.288744258652407e+17, 1.288744258693033e+17, 1.288744258732095e+17, 1.288744258772721e+17, 1.288744258813345e+17, 1.288744258852408e+17, 1.288744258893033e+17, 1.288744258932095e+17, 1.288744258972721e+17, 1.288744259013344e+17, 1.288744259052407e+17, 1.288744259093032e+17, 1.288744259132095e+17, 1.288744259172721e+17, 1.288744259213345e+17, 1.288744259252408e+17, 1.288744259293032e+17, 1.288744259332096e+17, 1.288744259372719e+17, 1.288744259413344e+17, 1.288744259452408e+17, 1.288744259493032e+17, 1.288744259532095e+17, 1.288744259572719e+17, 1.288744259613345e+17, 1.288744259652407e+17, 1.288744259693033e+17, 1.288744259732096e+17, 1.288744259772719e+17, 1.288744259813345e+17, 1.288744259852407e+17, 1.288744259893032e+17, 1.288744259932095e+17, 1.288744259972719e+17, 1.288744260013345e+17, 1.288744260052407e+17, 1.288744260093033e+17, 1.288744260132095e+17, 1.288744260172719e+17, 1.288744260213345e+17, 1.288744260252407e+17, 1.288744260293033e+17, 1.288744260332095e+17, 1.288744260372719e+17, 1.288744260413345e+17, 1.288744260452407e+17, 1.288744260493033e+17, 1.288744260532095e+17, 1.288744260572721e+17, 1.288744260613345e+17, 1.288744260652407e+17, 1.288744260693033e+17, 1.288744260732095e+17, 1.288744260772719e+17, 1.288744260813345e+17, 1.288744260852407e+17, 1.288744260893033e+17, 1.288744260932095e+17, 1.288744260972721e+17, 1.288744261013345e+17, 1.288744261052408e+17, 1.288744261093033e+17, 1.288744261132095e+17, 1.288744261172721e+17, 1.288744261213344e+17, 1.288744261252407e+17, 1.288744261293033e+17, 1.288744261332095e+17, 1.288744261372721e+17, 1.288744261413345e+17, 1.288744261452408e+17, 1.288744261493032e+17, 1.288744261532095e+17, 1.288744261572721e+17, 1.288744261613344e+17, 1.288744261652408e+17, 1.288744261693032e+17, 1.288744261732095e+17, 1.288744261772719e+17, 1.288744261813345e+17, 1.288744261852408e+17, 1.288744261893032e+17, 1.288744261932096e+17, 1.288744261972719e+17, 1.288744262013345e+17, 1.288744262052407e+17, 1.288744262093032e+17, 1.288744262132095e+17, 1.288744262172719e+17, 1.288744262213345e+17, 1.288744262252407e+17, 1.288744262293033e+17, 1.288744262332095e+17, 1.288744262372719e+17, 1.288744262413345e+17, 1.288744262452407e+17, 1.288744262493032e+17, 1.288744262532095e+17, 1.288744262572719e+17, 1.288744262613345e+17, 1.288744262652407e+17, 1.288744262693033e+17, 1.288744262732095e+17, 1.288744262772719e+17, 1.288744262813345e+17, 1.288744262852407e+17, 1.288744262893033e+17, 1.288744262932095e+17, 1.288744262972719e+17, 1.288744263013345e+17, 1.288744263052407e+17, 1.288744263093033e+17, 1.288744263132095e+17, 1.288744263172721e+17, 1.288744263213345e+17, 1.288744263252407e+17, 1.288744263293033e+17, 1.288744263332095e+17, 1.288744263372719e+17, 1.288744263413345e+17, 1.288744263452407e+17, 1.288744263493033e+17, 1.288744263532095e+17, 1.288744263572721e+17, 1.288744263613345e+17, 1.288744263652408e+17, 1.288744263693033e+17, 1.288744263732095e+17, 1.288744263772721e+17, 1.288744263813344e+17, 1.288744263852407e+17, 1.288744263893033e+17, 1.288744263932095e+17, 1.288744263972721e+17, 1.288744264013345e+17, 1.288744264052408e+17, 1.288744264093032e+17, 1.288744264132095e+17, 1.288744264172721e+17, 1.288744264213344e+17, 1.288744264252408e+17, 1.288744264293032e+17, 1.288744264332095e+17, 1.288744264372719e+17, 1.288744264413345e+17, 1.288744264452408e+17, 1.288744264493032e+17, 1.288744264532096e+17, 1.288744264572719e+17, 1.288744264613345e+17, 1.288744264652407e+17, 1.288744264693032e+17, 1.288744264732095e+17, 1.288744264772719e+17, 1.288744264813345e+17, 1.288744264852407e+17, 1.288744264893033e+17, 1.288744264932095e+17, 1.288744264972719e+17, 1.288744265013345e+17, 1.288744265052407e+17, 1.288744265093032e+17, 1.288744265132095e+17, 1.288744265172719e+17, 1.288744265213345e+17, 1.288744265252407e+17, 1.288744265293033e+17, 1.288744265332095e+17, 1.288744265372719e+17, 1.288744265413345e+17, 1.288744265452407e+17, 1.288744265493033e+17, 1.288744265532095e+17, 1.288744265572719e+17, 1.288744265613345e+17, 1.288744265652407e+17, 1.288744265693033e+17, 1.288744265732095e+17, 1.288744265772721e+17, 1.288744265813345e+17, 1.288744265852407e+17, 1.288744265893033e+17, 1.288744265932095e+17, 1.288744265972719e+17, 1.288744266013345e+17, 1.288744266052407e+17, 1.288744266093033e+17, 1.288744266132095e+17, 1.288744266172721e+17, 1.288744266213345e+17, 1.288744266252408e+17, 1.288744266293033e+17, 1.288744266332095e+17, 1.288744266372721e+17, 1.288744266413344e+17, 1.288744266452407e+17, 1.288744266493033e+17, 1.288744266532095e+17, 1.288744266572721e+17, 1.288744266613345e+17, 1.288744266652408e+17, 1.288744266693032e+17, 1.288744266732095e+17, 1.288744266772721e+17, 1.288744266813344e+17, 1.288744266852408e+17, 1.288744266893032e+17, 1.288744266932095e+17, 1.288744266972719e+17, 1.288744267013345e+17, 1.288744267052408e+17, 1.288744267093032e+17, 1.288744267132096e+17, 1.288744267172719e+17, 1.288744267213345e+17, 1.288744267252407e+17, 1.288744267293032e+17, 1.288744267332095e+17, 1.288744267372719e+17, 1.288744267413345e+17, 1.288744267452407e+17, 1.288744267493033e+17, 1.288744267532095e+17, 1.288744267572719e+17, 1.288744267613345e+17, 1.288744267652407e+17, 1.288744267693032e+17, 1.288744267732095e+17, 1.288744267772719e+17, 1.288744267813345e+17, 1.288744267852407e+17, 1.288744267893033e+17, 1.288744267932095e+17, 1.288744267972721e+17, 1.288744268013345e+17, 1.288744268052407e+17, 1.288744268093033e+17, 1.288744268132095e+17, 1.288744268172719e+17, 1.288744268213345e+17, 1.288744268252407e+17, 1.288744268293033e+17, 1.288744268332095e+17, 1.288744268372721e+17, 1.288744268413345e+17, 1.288744268452407e+17, 1.288744268493033e+17, 1.288744268532095e+17, 1.288744268572721e+17, 1.288744268613345e+17, 1.288744268652407e+17, 1.288744268693033e+17, 1.288744268732095e+17, 1.288744268772721e+17, 1.288744268813345e+17, 1.288744268852408e+17, 1.288744268893033e+17, 1.288744268932095e+17, 1.288744268972721e+17, 1.288744269013344e+17, 1.288744269052407e+17, 1.288744269093033e+17, 1.288744269132095e+17, 1.288744269172721e+17, 1.288744269213345e+17, 1.288744269252408e+17, 1.288744269293032e+17, 1.288744269332095e+17, 1.288744269372721e+17, 1.288744269413344e+17, 1.288744269452408e+17, 1.288744269493032e+17, 1.288744269532095e+17, 1.288744269572719e+17, 1.288744269613345e+17, 1.288744269652408e+17, 1.288744269693032e+17, 1.288744269732096e+17, 1.288744269772719e+17, 1.288744269813345e+17, 1.288744269852407e+17, 1.288744269893032e+17, 1.288744269932095e+17, 1.288744269972719e+17, 1.288744270013345e+17, 1.288744270052407e+17, 1.288744270093033e+17, 1.288744270132095e+17, 1.288744270172719e+17, 1.288744270213345e+17, 1.288744270252407e+17, 1.288744270293032e+17, 1.288744270332095e+17, 1.288744270372719e+17, 1.288744270413345e+17, 1.288744270452407e+17, 1.288744270493033e+17, 1.288744270532095e+17, 1.288744270572721e+17, 1.288744270613345e+17, 1.288744270652407e+17, 1.288744270693033e+17, 1.288744270732095e+17, 1.288744270772719e+17, 1.288744270813345e+17, 1.288744270852407e+17, 1.288744270893033e+17, 1.288744270932095e+17, 1.288744270972721e+17, 1.288744271013345e+17, 1.288744271052407e+17, 1.288744271093033e+17, 1.288744271132095e+17, 1.288744271172721e+17, 1.288744271213345e+17, 1.288744271252407e+17, 1.288744271293033e+17, 1.288744271332095e+17, 1.288744271372721e+17, 1.288744271413344e+17, 1.288744271452408e+17, 1.288744271493033e+17, 1.288744271532095e+17, 1.288744271572721e+17, 1.288744271613344e+17, 1.288744271652407e+17, 1.288744271693032e+17, 1.288744271732095e+17, 1.288744271772721e+17, 1.288744271813345e+17, 1.288744271852408e+17, 1.288744271893032e+17, 1.288744271932095e+17, 1.288744271972719e+17, 1.288744272013344e+17, 1.288744272052408e+17, 1.288744272093032e+17, 1.288744272132095e+17, 1.288744272172719e+17, 1.288744272213345e+17, 1.288744272252407e+17, 1.288744272293033e+17, 1.288744272332096e+17, 1.288744272372719e+17, 1.288744272413345e+17, 1.288744272452407e+17, 1.288744272493032e+17, 1.288744272532095e+17, 1.288744272572719e+17, 1.288744272613345e+17, 1.288744272652407e+17, 1.288744272693033e+17, 1.288744272732095e+17, 1.288744272772719e+17, 1.288744272813345e+17, 1.288744272852407e+17, 1.288744272893032e+17, 1.288744272932095e+17, 1.288744272972719e+17, 1.288744273013345e+17, 1.288744273052407e+17, 1.288744273093033e+17, 1.288744273132095e+17, 1.288744273172721e+17, 1.288744273213345e+17, 1.288744273252407e+17, 1.288744273293033e+17, 1.288744273332095e+17, 1.288744273372719e+17, 1.288744273413345e+17, 1.288744273452407e+17, 1.288744273493033e+17, 1.288744273532095e+17, 1.288744273572721e+17, 1.288744273613345e+17, 1.288744273652407e+17, 1.288744273693033e+17, 1.288744273732095e+17, 1.288744273772721e+17, 1.288744273813345e+17, 1.288744273852407e+17, 1.288744273893033e+17, 1.288744273932095e+17, 1.288744273972721e+17, 1.288744274013344e+17, 1.288744274052408e+17, 1.288744274093033e+17, 1.288744274132095e+17, 1.288744274172721e+17, 1.288744274213344e+17, 1.288744274252407e+17, 1.288744274293032e+17, 1.288744274332095e+17, 1.288744274372721e+17, 1.288744274413345e+17, 1.288744274452408e+17, 1.288744274493032e+17, 1.288744274532096e+17, 1.288744274572719e+17, 1.288744274613344e+17, 1.288744274652408e+17, 1.288744274693032e+17, 1.288744274732095e+17, 1.288744274772719e+17, 1.288744274813345e+17, 1.288744274852407e+17, 1.288744274893033e+17, 1.288744274932096e+17, 1.288744274972719e+17, 1.288744275013345e+17, 1.288744275052407e+17, 1.288744275093032e+17, 1.288744275132095e+17, 1.288744275172719e+17, 1.288744275213345e+17, 1.288744275252407e+17, 1.288744275293033e+17, 1.288744275332095e+17, 1.288744275372719e+17, 1.288744275413345e+17, 1.288744275452407e+17, 1.288744275493033e+17, 1.288744275532095e+17, 1.288744275572719e+17, 1.288744275613345e+17, 1.288744275652407e+17, 1.288744275693033e+17, 1.288744275732095e+17, 1.288744275772721e+17, 1.288744275813345e+17, 1.288744275852407e+17, 1.288744275893033e+17, 1.288744275932095e+17, 1.288744275972719e+17, 1.288744276013345e+17, 1.288744276052407e+17, 1.288744276093033e+17, 1.288744276132095e+17, 1.288744276172721e+17, 1.288744276213345e+17, 1.288744276252407e+17, 1.288744276293033e+17, 1.288744276332095e+17, 1.288744276372721e+17, 1.288744276413345e+17, 1.288744276452407e+17, 1.288744276493033e+17, 1.288744276532095e+17, 1.288744276572721e+17, 1.288744276613344e+17, 1.288744276652408e+17, 1.288744276693033e+17, 1.288744276732095e+17, 1.288744276772721e+17, 1.288744276813344e+17, 1.288744276852407e+17, 1.288744276893032e+17, 1.288744276932095e+17, 1.288744276972721e+17, 1.288744277013345e+17, 1.288744277052408e+17, 1.288744277093032e+17, 1.288744277132096e+17, 1.288744277172719e+17, 1.288744277213344e+17, 1.288744277252408e+17, 1.288744277293032e+17, 1.288744277332095e+17, 1.288744277372719e+17, 1.288744277413345e+17, 1.288744277452407e+17, 1.288744277493033e+17, 1.288744277532096e+17, 1.288744277572719e+17, 1.288744277613345e+17, 1.288744277652407e+17, 1.288744277693032e+17, 1.288744277732095e+17, 1.288744277772719e+17, 1.288744277813345e+17, 1.288744277852407e+17, 1.288744277893033e+17, 1.288744277932095e+17, 1.288744277972719e+17, 1.288744278013345e+17, 1.288744278052407e+17, 1.288744278093033e+17, 1.288744278132095e+17, 1.288744278172719e+17, 1.288744278213345e+17, 1.288744278252407e+17, 1.288744278293033e+17, 1.288744278332095e+17, 1.288744278372721e+17, 1.288744278413345e+17, 1.288744278452407e+17, 1.288744278493033e+17, 1.288744278532095e+17, 1.288744278572719e+17, 1.288744278613345e+17, 1.288744278652407e+17, 1.288744278693033e+17, 1.288744278732095e+17, 1.288744278772721e+17, 1.288744278813345e+17, 1.288744278852408e+17, 1.288744278893033e+17, 1.288744278932095e+17, 1.288744278972721e+17, 1.288744279013345e+17, 1.288744279052407e+17, 1.288744279093033e+17, 1.288744279132095e+17, 1.288744279172721e+17, 1.288744279213345e+17, 1.288744279252408e+17, 1.288744279293033e+17, 1.288744279332095e+17, 1.288744279372721e+17, 1.288744279413344e+17, 1.288744279452407e+17, 1.288744279493032e+17, 1.288744279532095e+17, 1.288744279572721e+17, 1.288744279613345e+17, 1.288744279652408e+17, 1.288744279693032e+17, 1.288744279732096e+17, 1.288744279772719e+17, 1.288744279813344e+17, 1.288744279852408e+17, 1.288744279893032e+17, 1.288744279932095e+17, 1.288744279972719e+17, 1.288744280013345e+17, 1.288744280052407e+17, 1.288744280093033e+17, 1.288744280132096e+17, 1.288744280172719e+17, 1.288744280213345e+17, 1.288744280252407e+17, 1.288744280293032e+17, 1.288744280332095e+17, 1.288744280372719e+17, 1.288744280413345e+17, 1.288744280452407e+17, 1.288744280493033e+17, 1.288744280532095e+17, 1.288744280572719e+17, 1.288744280613345e+17, 1.288744280652407e+17, 1.288744280693033e+17, 1.288744280732095e+17, 1.288744280772719e+17, 1.288744280813345e+17, 1.288744280852407e+17, 1.288744280893033e+17, 1.288744280932095e+17, 1.288744280972721e+17, 1.288744281013345e+17, 1.288744281052407e+17, 1.288744281093033e+17, 1.288744281132095e+17, 1.288744281172719e+17, 1.288744281213345e+17, 1.288744281252407e+17, 1.288744281293033e+17, 1.288744281332095e+17, 1.288744281372721e+17, 1.288744281413345e+17, 1.288744281452408e+17, 1.288744281493033e+17, 1.288744281532095e+17, 1.288744281572721e+17, 1.288744281613344e+17, 1.288744281652407e+17, 1.288744281693033e+17, 1.288744281732095e+17, 1.288744281772721e+17, 1.288744281813345e+17, 1.288744281852408e+17, 1.288744281893032e+17, 1.288744281932095e+17, 1.288744281972721e+17, 1.288744282013344e+17, 1.288744282052408e+17, 1.288744282093032e+17, 1.288744282132095e+17, 1.288744282172719e+17, 1.288744282213345e+17, 1.288744282252408e+17, 1.288744282293032e+17, 1.288744282332096e+17, 1.288744282372719e+17, 1.288744282413345e+17, 1.288744282452407e+17, 1.288744282493032e+17, 1.288744282532095e+17, 1.288744282572719e+17, 1.288744282613345e+17, 1.288744282652407e+17, 1.288744282693033e+17, 1.288744282732095e+17, 1.288744282772719e+17, 1.288744282813345e+17, 1.288744282852407e+17, 1.288744282893032e+17, 1.288744282932095e+17, 1.288744282972719e+17, 1.288744283013345e+17, 1.288744283052407e+17, 1.288744283093033e+17, 1.288744283132095e+17, 1.288744283172719e+17, 1.288744283213345e+17, 1.288744283252407e+17, 1.288744283293033e+17, 1.288744283332095e+17, 1.288744283372719e+17, 1.288744283413345e+17, 1.288744283452407e+17, 1.288744283493033e+17, 1.288744283532095e+17, 1.288744283572721e+17, 1.288744283613345e+17, 1.288744283652407e+17, 1.288744283693033e+17, 1.288744283732095e+17, 1.288744283772719e+17, 1.288744283813345e+17, 1.288744283852407e+17, 1.288744283893033e+17, 1.288744283932095e+17, 1.288744283972721e+17, 1.288744284013345e+17, 1.288744284052408e+17, 1.288744284093033e+17, 1.288744284132095e+17, 1.288744284172721e+17, 1.288744284213344e+17, 1.288744284252407e+17, 1.288744284293033e+17, 1.288744284332095e+17, 1.288744284372721e+17, 1.288744284413345e+17, 1.288744284452408e+17, 1.288744284493032e+17, 1.288744284532095e+17, 1.288744284572721e+17, 1.288744284613344e+17, 1.288744284652408e+17, 1.288744284693032e+17, 1.288744284732095e+17, 1.288744284772719e+17, 1.288744284813345e+17, 1.288744284852408e+17, 1.288744284893032e+17, 1.288744284932096e+17, 1.288744284972719e+17, 1.288744285013345e+17, 1.288744285052407e+17, 1.288744285093032e+17, 1.288744285132095e+17, 1.288744285172719e+17, 1.288744285213345e+17, 1.288744285252407e+17, 1.288744285293033e+17, 1.288744285332095e+17, 1.288744285372719e+17, 1.288744285413345e+17, 1.288744285452407e+17, 1.288744285493032e+17, 1.288744285532095e+17, 1.288744285572719e+17, 1.288744285613345e+17, 1.288744285652407e+17, 1.288744285693033e+17, 1.288744285732095e+17, 1.288744285772721e+17, 1.288744285813345e+17, 1.288744285852407e+17, 1.288744285893033e+17, 1.288744285932095e+17, 1.288744285972719e+17, 1.288744286013345e+17, 1.288744286052407e+17, 1.288744286093033e+17, 1.288744286132095e+17, 1.288744286172721e+17, 1.288744286213345e+17, 1.288744286252407e+17, 1.288744286293033e+17, 1.288744286332095e+17, 1.288744286372719e+17, 1.288744286413345e+17, 1.288744286452407e+17, 1.288744286493033e+17, 1.288744286532095e+17, 1.288744286572721e+17, 1.288744286613345e+17, 1.288744286652408e+17, 1.288744286693033e+17, 1.288744286732095e+17, 1.288744286772721e+17, 1.288744286813344e+17, 1.288744286852407e+17, 1.288744286893033e+17, 1.288744286932095e+17, 1.288744286972721e+17, 1.288744287013345e+17, 1.288744287052408e+17, 1.288744287093032e+17, 1.288744287132095e+17, 1.288744287172721e+17, 1.288744287213344e+17, 1.288744287252408e+17, 1.288744287293032e+17, 1.288744287332095e+17, 1.288744287372719e+17, 1.288744287413345e+17, 1.288744287452408e+17, 1.288744287493032e+17, 1.288744287532096e+17, 1.288744287572719e+17, 1.288744287613345e+17, 1.288744287652407e+17, 1.288744287693032e+17, 1.288744287732095e+17, 1.288744287772719e+17, 1.288744287813345e+17, 1.288744287852407e+17, 1.288744287893033e+17, 1.288744287932095e+17, 1.288744287972719e+17, 1.288744288013345e+17, 1.288744288052407e+17, 1.288744288093032e+17, 1.288744288132095e+17, 1.288744288172719e+17, 1.288744288213345e+17, 1.288744288252407e+17, 1.288744288293033e+17, 1.288744288332095e+17, 1.288744288372721e+17, 1.288744288413345e+17, 1.288744288452407e+17, 1.288744288493033e+17, 1.288744288532095e+17, 1.288744288572719e+17, 1.288744288613345e+17, 1.288744288652407e+17, 1.288744288693033e+17, 1.288744288732095e+17, 1.288744288772721e+17, 1.288744288813345e+17, 1.288744288852407e+17, 1.288744288893033e+17, 1.288744288932095e+17, 1.288744288972721e+17, 1.288744289013345e+17, 1.288744289052407e+17, 1.288744289093033e+17, 1.288744289132095e+17, 1.288744289172721e+17, 1.288744289213345e+17, 1.288744289252408e+17, 1.288744289293033e+17, 1.288744289332095e+17, 1.288744289372721e+17, 1.288744289413344e+17, 1.288744289452407e+17, 1.288744289493033e+17, 1.288744289532095e+17, 1.288744289572721e+17, 1.288744289613345e+17, 1.288744289652408e+17, 1.288744289693032e+17, 1.288744289732095e+17, 1.288744289772721e+17, 1.288744289813344e+17, 1.288744289852408e+17, 1.288744289893032e+17, 1.288744289932095e+17, 1.288744289972719e+17, 1.288744290013345e+17, 1.288744290052408e+17, 1.288744290093032e+17, 1.288744290132096e+17, 1.288744290172719e+17, 1.288744290213345e+17, 1.288744290252407e+17, 1.288744290293032e+17, 1.288744290332095e+17, 1.288744290372719e+17, 1.288744290413345e+17, 1.288744290452407e+17, 1.288744290493033e+17, 1.288744290532095e+17, 1.288744290572719e+17, 1.288744290613345e+17, 1.288744290652407e+17, 1.288744290693032e+17, 1.288744290732095e+17, 1.288744290772719e+17, 1.288744290813345e+17, 1.288744290852407e+17, 1.288744290893033e+17, 1.288744290932095e+17, 1.288744290972721e+17, 1.288744291013345e+17, 1.288744291052407e+17, 1.288744291093033e+17, 1.288744291132095e+17, 1.288744291172719e+17, 1.288744291213345e+17, 1.288744291252407e+17, 1.288744291293033e+17, 1.288744291332095e+17, 1.288744291372721e+17, 1.288744291413345e+17, 1.288744291452407e+17, 1.288744291493033e+17, 1.288744291532095e+17, 1.288744291572721e+17, 1.288744291613345e+17, 1.288744291652407e+17, 1.288744291693033e+17, 1.288744291732095e+17, 1.288744291772721e+17, 1.288744291813344e+17, 1.288744291852408e+17, 1.288744291893033e+17, 1.288744291932095e+17, 1.288744291972721e+17, 1.288744292013344e+17, 1.288744292052407e+17, 1.288744292093032e+17, 1.288744292132095e+17, 1.288744292172721e+17, 1.288744292213345e+17, 1.288744292252408e+17, 1.288744292293032e+17, 1.288744292332096e+17, 1.288744292372719e+17, 1.288744292413344e+17, 1.288744292452408e+17, 1.288744292493032e+17, 1.288744292532095e+17, 1.288744292572719e+17, 1.288744292613345e+17, 1.288744292652407e+17, 1.288744292693033e+17, 1.288744292732096e+17, 1.288744292772719e+17, 1.288744292813345e+17, 1.288744292852407e+17, 1.288744292893032e+17, 1.288744292932095e+17, 1.288744292972719e+17, 1.288744293013345e+17, 1.288744293052407e+17, 1.288744293093033e+17, 1.288744293132095e+17, 1.288744293172719e+17, 1.288744293213345e+17, 1.288744293252407e+17, 1.288744293293033e+17, 1.288744293332095e+17, 1.288744293372719e+17, 1.288744293413345e+17, 1.288744293452407e+17, 1.288744293493033e+17, 1.288744293532095e+17, 1.288744293572721e+17, 1.288744293613345e+17, 1.288744293652407e+17, 1.288744293693033e+17, 1.288744293732095e+17, 1.288744293772719e+17, 1.288744293813345e+17, 1.288744293852407e+17, 1.288744293893033e+17, 1.288744293932095e+17, 1.288744293972721e+17, 1.288744294013345e+17, 1.288744294052407e+17, 1.288744294093033e+17, 1.288744294132095e+17, 1.288744294172721e+17, 1.288744294213345e+17, 1.288744294252407e+17, 1.288744294293033e+17, 1.288744294413344e+17, 1.288744294452408e+17, 1.288744294493033e+17, 1.288744294532095e+17, 1.288744294572721e+17, 1.288744294613344e+17, 1.288744294652407e+17, 1.288744294693032e+17, 1.288744294732095e+17, 1.288744294772721e+17, 1.288744294813345e+17, 1.288744294852408e+17, 1.288744294893032e+17, 1.288744294932096e+17, 1.288744294972719e+17, 1.288744295013344e+17, 1.288744295052408e+17, 1.288744295093032e+17, 1.288744295132095e+17, 1.288744295172719e+17, 1.288744295213345e+17, 1.288744295252407e+17, 1.288744295293033e+17, 1.288744295332096e+17, 1.288744295372719e+17, 1.288744295413345e+17, 1.288744295452407e+17, 1.288744295493032e+17, 1.288744295532095e+17, 1.288744295572719e+17, 1.288744295613345e+17, 1.288744295652407e+17, 1.288744295693033e+17, 1.288744295732095e+17, 1.288744295772719e+17, 1.288744295813345e+17, 1.288744295852407e+17, 1.288744295893033e+17, 1.288744295932095e+17, 1.288744295972719e+17, 1.288744296013345e+17, 1.288744296052407e+17, 1.288744296093033e+17, 1.288744296132095e+17, 1.288744296172721e+17, 1.288744296213345e+17, 1.288744296252407e+17, 1.288744296293033e+17, 1.288744296332095e+17, 1.288744296372719e+17, 1.288744296413345e+17, 1.288744296452407e+17, 1.288744296493033e+17, 1.288744296532095e+17, 1.288744296572721e+17, 1.288744296613345e+17, 1.288744296652407e+17, 1.288744296693033e+17, 1.288744296732095e+17, 1.288744296772721e+17, 1.288744296813345e+17, 1.288744296852407e+17, 1.288744296893033e+17, 1.288744296932095e+17, 1.288744296972721e+17, 1.288744297013344e+17, 1.288744297052408e+17, 1.288744297093033e+17, 1.288744297132095e+17, 1.288744297172721e+17, 1.288744297213344e+17, 1.288744297252407e+17, 1.288744297293032e+17, 1.288744297332095e+17, 1.288744297372721e+17, 1.288744297413345e+17, 1.288744297452408e+17, 1.288744297493032e+17, 1.288744297532096e+17, 1.288744297572719e+17, 1.288744297613344e+17, 1.288744297652408e+17, 1.288744297693032e+17, 1.288744297732095e+17, 1.288744297772719e+17, 1.288744297813345e+17, 1.288744297852407e+17, 1.288744297893033e+17, 1.288744297932096e+17, 1.288744297972719e+17, 1.288744298013345e+17, 1.288744298052407e+17, 1.288744298093032e+17, 1.288744298132095e+17, 1.288744298172719e+17, 1.288744298213345e+17, 1.288744298252407e+17, 1.288744298293033e+17, 1.288744298332095e+17, 1.288744298372719e+17, 1.288744298413345e+17, 1.288744298452407e+17, 1.288744298493033e+17, 1.288744298532095e+17, 1.288744298572719e+17, 1.288744298613345e+17, 1.288744298652407e+17, 1.288744298693033e+17, 1.288744298732095e+17, 1.288744298772721e+17, 1.288744298813345e+17, 1.288744298852407e+17, 1.288744298893033e+17, 1.288744298932095e+17, 1.288744298972719e+17, 1.288744299013345e+17, 1.288744299052407e+17, 1.288744299093033e+17, 1.288744299132095e+17, 1.288744299172721e+17, 1.288744299213345e+17, 1.288744299252408e+17, 1.288744299293033e+17, 1.288744299332095e+17, 1.288744299372721e+17, 1.288744299413344e+17, 1.288744299452407e+17, 1.288744299493033e+17, 1.288744299532095e+17, 1.288744299572721e+17, 1.288744299613345e+17, 1.288744299652408e+17, 1.288744299693032e+17, 1.288744299732095e+17, 1.288744299772721e+17, 1.288744299813344e+17, 1.288744299852407e+17, 1.288744299893032e+17, 1.288744299932095e+17, 1.288744299972719e+17, 1.288744300013345e+17, 1.288744300052408e+17, 1.288744300093032e+17, 1.288744300132096e+17, 1.288744300172719e+17, 1.288744300213345e+17, 1.288744300252407e+17, 1.288744300293032e+17, 1.288744300332095e+17, 1.288744300372719e+17, 1.288744300413345e+17, 1.288744300452407e+17, 1.288744300493033e+17, 1.288744300532095e+17, 1.288744300572719e+17, 1.288744300613345e+17, 1.288744300652407e+17, 1.288744300693032e+17, 1.288744300732095e+17, 1.288744300772719e+17, 1.288744300813345e+17, 1.288744300852407e+17, 1.288744300893033e+17, 1.288744300932095e+17, 1.288744300972719e+17, 1.288744301013345e+17, 1.288744301052407e+17, 1.288744301093033e+17, 1.288744301132095e+17, 1.288744301172719e+17, 1.288744301213345e+17, 1.288744301252407e+17, 1.288744301293033e+17, 1.288744301332095e+17, 1.288744301372721e+17, 1.288744301413345e+17, 1.288744301452407e+17, 1.288744301493033e+17, 1.288744301532095e+17, 1.288744301572719e+17, 1.288744301613345e+17, 1.288744301652407e+17, 1.288744301693033e+17, 1.288744301732095e+17, 1.288744301772721e+17, 1.288744301813345e+17, 1.288744301852408e+17, 1.288744301893033e+17, 1.288744301932095e+17, 1.288744301972721e+17, 1.288744302013344e+17, 1.288744302052407e+17, 1.288744302093033e+17, 1.288744302132095e+17, 1.288744302172721e+17, 1.288744302213345e+17, 1.288744302252408e+17, 1.288744302293032e+17, 1.288744302332095e+17, 1.288744302372721e+17, 1.288744302413344e+17, 1.288744302452408e+17, 1.288744302493032e+17, 1.288744302532095e+17, 1.288744302572719e+17, 1.288744302613345e+17, 1.288744302652408e+17, 1.288744302693032e+17, 1.288744302732096e+17, 1.288744302772719e+17, 1.288744302813345e+17, 1.288744302852407e+17, 1.288744302893032e+17, 1.288744302932095e+17, 1.288744302972719e+17, 1.288744303013345e+17, 1.288744303052407e+17, 1.288744303093033e+17, 1.288744303132095e+17, 1.288744303172719e+17, 1.288744303213345e+17, 1.288744303252407e+17, 1.288744303293032e+17, 1.288744303332095e+17, 1.288744303372719e+17, 1.288744303413345e+17, 1.288744303452407e+17, 1.288744303493033e+17, 1.288744303532095e+17, 1.288744303572719e+17, 1.288744303613345e+17, 1.288744303652407e+17, 1.288744303693033e+17, 1.288744303732095e+17, 1.288744303772719e+17, 1.288744303813345e+17, 1.288744303852407e+17, 1.288744303893033e+17, 1.288744303932095e+17, 1.288744303972721e+17, 1.288744304013345e+17, 1.288744304052407e+17, 1.288744304093033e+17, 1.288744304132095e+17, 1.288744304172719e+17, 1.288744304213345e+17, 1.288744304252407e+17, 1.288744304293033e+17, 1.288744304332095e+17, 1.288744304372721e+17, 1.288744304413345e+17, 1.288744304452408e+17, 1.288744304493033e+17, 1.288744304532095e+17, 1.288744304572721e+17, 1.288744304613344e+17, 1.288744304652407e+17, 1.288744304693033e+17, 1.288744304732095e+17, 1.288744304772721e+17, 1.288744304813345e+17, 1.288744304852408e+17, 1.288744304893032e+17, 1.288744304932095e+17, 1.288744304972721e+17, 1.288744305013344e+17, 1.288744305052408e+17, 1.288744305093032e+17, 1.288744305132095e+17, 1.288744305172719e+17, 1.288744305213345e+17, 1.288744305252408e+17, 1.288744305293032e+17, 1.288744305332096e+17, 1.288744305372719e+17, 1.288744305413345e+17, 1.288744305452407e+17, 1.288744305493032e+17, 1.288744305532095e+17, 1.288744305572719e+17, 1.288744305613345e+17, 1.288744305652407e+17, 1.288744305693033e+17, 1.288744305732095e+17, 1.288744305772719e+17, 1.288744305813345e+17, 1.288744305852407e+17, 1.288744305893032e+17, 1.288744305932095e+17, 1.288744305972719e+17, 1.288744306013345e+17, 1.288744306052407e+17, 1.288744306093033e+17, 1.288744306132095e+17, 1.288744306172721e+17, 1.288744306213345e+17, 1.288744306252407e+17, 1.288744306293033e+17, 1.288744306332095e+17, 1.288744306372719e+17, 1.288744306413345e+17, 1.288744306452407e+17, 1.288744306493033e+17, 1.288744306532095e+17, 1.288744306572721e+17, 1.288744306613345e+17, 1.288744306652407e+17, 1.288744306693033e+17, 1.288744306732095e+17, 1.288744306772721e+17, 1.288744306813345e+17, 1.288744306852407e+17, 1.288744306893033e+17, 1.288744306932095e+17, 1.288744306972721e+17, 1.288744307013345e+17, 1.288744307052408e+17, 1.288744307093033e+17, 1.288744307132095e+17, 1.288744307172721e+17, 1.288744307213344e+17, 1.288744307252407e+17, 1.288744307293033e+17, 1.288744307332095e+17, 1.288744307372721e+17, 1.288744307413345e+17, 1.288744307452408e+17, 1.288744307493032e+17, 1.288744307532095e+17, 1.288744307572721e+17, 1.288744307613344e+17, 1.288744307652408e+17, 1.288744307693032e+17, 1.288744307732095e+17, 1.288744307772719e+17, 1.288744307813345e+17, 1.288744307852408e+17, 1.288744307893032e+17, 1.288744307932096e+17, 1.288744307972719e+17, 1.288744308013345e+17, 1.288744308052407e+17, 1.288744308093032e+17, 1.288744308132095e+17, 1.288744308172719e+17, 1.288744308213345e+17, 1.288744308252407e+17, 1.288744308293033e+17, 1.288744308332095e+17, 1.288744308372719e+17, 1.288744308413345e+17, 1.288744308452407e+17, 1.288744308493032e+17, 1.288744308532095e+17, 1.288744308572719e+17, 1.288744308613345e+17, 1.288744308652407e+17, 1.288744308693033e+17, 1.288744308732095e+17, 1.288744308772721e+17, 1.288744308813345e+17, 1.288744308852407e+17, 1.288744308893033e+17, 1.288744308932095e+17, 1.288744308972719e+17, 1.288744309013345e+17, 1.288744309052407e+17, 1.288744309093033e+17, 1.288744309132095e+17, 1.288744309172721e+17, 1.288744309213345e+17, 1.288744309252407e+17, 1.288744309293033e+17, 1.288744309332095e+17, 1.288744309372721e+17, 1.288744309413345e+17, 1.288744309452407e+17, 1.288744309493033e+17, 1.288744309532095e+17, 1.288744309572721e+17, 1.288744309613344e+17, 1.288744309652408e+17, 1.288744309693033e+17, 1.288744309732095e+17, 1.288744309772721e+17, 1.288744309813344e+17, 1.288744309852407e+17, 1.288744309893032e+17, 1.288744309932095e+17, 1.288744309972721e+17, 1.288744310013345e+17, 1.288744310052408e+17, 1.288744310093032e+17, 1.288744310132095e+17, 1.288744310172719e+17, 1.288744310213344e+17, 1.288744310252408e+17, 1.288744310293032e+17, 1.288744310332095e+17, 1.288744310372719e+17, 1.288744310413345e+17, 1.288744310452407e+17, 1.288744310493033e+17, 1.288744310532096e+17, 1.288744310572719e+17, 1.288744310613345e+17, 1.288744310652407e+17, 1.288744310693032e+17, 1.288744310732095e+17, 1.288744310772719e+17, 1.288744310813345e+17, 1.288744310852407e+17, 1.288744310893033e+17, 1.288744310932095e+17, 1.288744310972719e+17, 1.288744311013345e+17, 1.288744311052407e+17, 1.288744311093032e+17, 1.288744311132095e+17, 1.288744311172719e+17, 1.288744311213345e+17, 1.288744311252407e+17, 1.288744311293033e+17, 1.288744311332095e+17, 1.288744311372721e+17, 1.288744311413345e+17, 1.288744311452407e+17, 1.288744311493033e+17, 1.288744311532095e+17, 1.288744311572719e+17, 1.288744311613345e+17, 1.288744311652407e+17, 1.288744311693033e+17, 1.288744311732095e+17, 1.288744311772721e+17, 1.288744311813345e+17, 1.288744311852407e+17, 1.288744311893033e+17, 1.288744311932095e+17, 1.288744311972721e+17, 1.288744312013345e+17, 1.288744312052407e+17, 1.288744312093033e+17, 1.288744312132095e+17, 1.288744312172721e+17, 1.288744312213344e+17, 1.288744312252408e+17, 1.288744312293033e+17, 1.288744312332095e+17, 1.288744312372721e+17, 1.288744312413344e+17, 1.288744312452407e+17, 1.288744312493032e+17, 1.288744312532095e+17, 1.288744312572721e+17, 1.288744312613345e+17, 1.288744312652408e+17, 1.288744312693032e+17, 1.288744312732096e+17, 1.288744312772719e+17, 1.288744312813344e+17, 1.288744312852408e+17, 1.288744312893032e+17, 1.288744312932095e+17, 1.288744312972719e+17, 1.288744313013345e+17, 1.288744313052407e+17, 1.288744313093033e+17, 1.288744313132096e+17, 1.288744313172719e+17, 1.288744313213345e+17, 1.288744313252407e+17, 1.288744313293032e+17, 1.288744313332095e+17, 1.288744313372719e+17, 1.288744313413345e+17, 1.288744313452407e+17, 1.288744313493033e+17, 1.288744313532095e+17, 1.288744313572719e+17, 1.288744313613345e+17, 1.288744313652407e+17, 1.288744313693033e+17, 1.288744313732095e+17, 1.288744313772719e+17, 1.288744313813345e+17, 1.288744313852407e+17, 1.288744313893033e+17, 1.288744313932095e+17, 1.288744313972721e+17, 1.288744314013345e+17, 1.288744314052407e+17, 1.288744314093033e+17, 1.288744314132095e+17, 1.288744314172719e+17, 1.288744314213345e+17, 1.288744314252407e+17, 1.288744314293033e+17, 1.288744314332095e+17, 1.288744314372721e+17, 1.288744314413345e+17, 1.288744314452407e+17, 1.288744314493033e+17, 1.288744314532095e+17, 1.288744314572721e+17, 1.288744314613345e+17, 1.288744314652407e+17, 1.288744314693033e+17, 1.288744314732095e+17, 1.288744314772721e+17, 1.288744314813344e+17, 1.288744314852408e+17, 1.288744314893033e+17, 1.288744314932095e+17, 1.288744314972721e+17, 1.288744315013344e+17, 1.288744315052407e+17, 1.288744315093032e+17, 1.288744315132095e+17, 1.288744315172721e+17, 1.288744315213345e+17, 1.288744315252408e+17, 1.288744315293032e+17, 1.288744315332096e+17, 1.288744315372719e+17, 1.288744315413344e+17, 1.288744315452408e+17, 1.288744315493032e+17, 1.288744315532095e+17, 1.288744315572719e+17, 1.288744315613345e+17, 1.288744315652407e+17, 1.288744315693033e+17, 1.288744315732096e+17, 1.288744315772719e+17, 1.288744315813345e+17, 1.288744315852407e+17, 1.288744315893032e+17, 1.288744315932095e+17, 1.288744315972719e+17, 1.288744316013345e+17, 1.288744316052407e+17, 1.288744316093033e+17, 1.288744316132095e+17, 1.288744316172719e+17, 1.288744316213345e+17, 1.288744316252407e+17, 1.288744316293033e+17, 1.288744316332095e+17, 1.288744316372719e+17, 1.288744316413345e+17, 1.288744316452407e+17, 1.288744316493033e+17, 1.288744316532095e+17, 1.288744316572721e+17, 1.288744316613345e+17, 1.288744316652407e+17, 1.288744316693033e+17, 1.288744316732095e+17, 1.288744316772719e+17, 1.288744316813345e+17, 1.288744316852407e+17, 1.288744316893033e+17, 1.288744316932095e+17, 1.288744316972721e+17, 1.288744317013345e+17, 1.288744317052407e+17, 1.288744317093033e+17, 1.288744317132095e+17, 1.288744317172721e+17, 1.288744317213345e+17, 1.288744317252407e+17, 1.288744317293033e+17, 1.288744317332095e+17, 1.288744317372721e+17, 1.288744317413345e+17, 1.288744317452408e+17, 1.288744317493033e+17, 1.288744317532095e+17, 1.288744317572721e+17, 1.288744317613344e+17, 1.288744317652407e+17, 1.288744317693032e+17, 1.288744317732095e+17, 1.288744317772721e+17, 1.288744317813345e+17, 1.288744317852408e+17, 1.288744317893032e+17, 1.288744317932096e+17, 1.288744317972719e+17, 1.288744318013344e+17, 1.288744318052408e+17, 1.288744318093032e+17, 1.288744318132095e+17, 1.288744318172719e+17, 1.288744318213345e+17, 1.288744318252407e+17, 1.288744318293033e+17, 1.288744318332096e+17, 1.288744318372719e+17, 1.288744318413345e+17, 1.288744318452407e+17, 1.288744318493032e+17, 1.288744318532095e+17, 1.288744318572719e+17, 1.288744318613345e+17, 1.288744318652407e+17, 1.288744318693033e+17, 1.288744318732095e+17, 1.288744318772719e+17, 1.288744318813345e+17, 1.288744318852407e+17, 1.288744318893033e+17, 1.288744318932095e+17, 1.288744318972719e+17, 1.288744319013345e+17, 1.288744319052407e+17, 1.288744319093033e+17, 1.288744319132095e+17, 1.288744319172721e+17, 1.288744319213345e+17, 1.288744319252407e+17, 1.288744319293033e+17, 1.288744319332095e+17, 1.288744319372719e+17, 1.288744319413345e+17, 1.288744319452407e+17, 1.288744319493033e+17, 1.288744319532095e+17, 1.288744319572721e+17, 1.288744319613345e+17, 1.288744319652408e+17, 1.288744319693033e+17, 1.288744319732095e+17, 1.288744319772721e+17, 1.288744319813344e+17, 1.288744319852407e+17, 1.288744319893033e+17, 1.288744319932095e+17, 1.288744319972721e+17, 1.288744320013345e+17, 1.288744320052408e+17, 1.288744320093032e+17, 1.288744320132095e+17, 1.288744320172721e+17, 1.288744320213344e+17, 1.288744320252408e+17, 1.288744320293032e+17, 1.288744320332095e+17, 1.288744320372719e+17, 1.288744320413345e+17, 1.288744320452408e+17, 1.288744320493032e+17, 1.288744320532096e+17, 1.288744320572719e+17, 1.288744320613345e+17, 1.288744320652407e+17, 1.288744320693032e+17, 1.288744320732095e+17, 1.288744320772719e+17, 1.288744320813345e+17, 1.288744320852407e+17, 1.288744320893033e+17, 1.288744320932095e+17, 1.288744320972719e+17, 1.288744321013345e+17, 1.288744321052407e+17, 1.288744321093032e+17, 1.288744321132095e+17, 1.288744321172719e+17, 1.288744321213345e+17, 1.288744321252407e+17, 1.288744321293033e+17, 1.288744321332095e+17, 1.288744321372719e+17, 1.288744321413345e+17, 1.288744321452407e+17, 1.288744321493033e+17, 1.288744321532095e+17, 1.288744321572719e+17, 1.288744321613345e+17, 1.288744321652407e+17, 1.288744321693033e+17, 1.288744321732095e+17, 1.288744321772721e+17, 1.288744321813345e+17, 1.288744321852407e+17, 1.288744321893033e+17, 1.288744321932095e+17, 1.288744321972719e+17, 1.288744322013345e+17, 1.288744322052407e+17, 1.288744322093033e+17, 1.288744322132095e+17, 1.288744322172721e+17, 1.288744322213345e+17, 1.288744322252408e+17, 1.288744322293033e+17, 1.288744322332095e+17, 1.288744322372721e+17, 1.288744322413344e+17, 1.288744322452407e+17, 1.288744322493033e+17, 1.288744322532095e+17, 1.288744322572721e+17, 1.288744322613345e+17, 1.288744322652408e+17, 1.288744322693032e+17, 1.288744322732095e+17, 1.288744322772721e+17, 1.288744322813344e+17, 1.288744322852408e+17, 1.288744322893032e+17, 1.288744322932095e+17, 1.288744322972719e+17, 1.288744323013345e+17, 1.288744323052408e+17, 1.288744323093032e+17, 1.288744323132096e+17, 1.288744323172719e+17, 1.288744323213345e+17, 1.288744323252407e+17, 1.288744323293032e+17, 1.288744323332095e+17, 1.288744323372719e+17, 1.288744323413345e+17, 1.288744323452407e+17, 1.288744323493033e+17, 1.288744323532095e+17, 1.288744323572719e+17, 1.288744323613345e+17, 1.288744323652407e+17, 1.288744323693032e+17, 1.288744323732095e+17, 1.288744323772719e+17, 1.288744323813345e+17, 1.288744323852407e+17, 1.288744323893033e+17, 1.288744323932095e+17, 1.288744323972721e+17, 1.288744324013345e+17, 1.288744324052407e+17, 1.288744324093033e+17, 1.288744324132095e+17, 1.288744324172719e+17, 1.288744324213345e+17, 1.288744324252407e+17, 1.288744324293033e+17, 1.288744324332095e+17, 1.288744324372721e+17, 1.288744324413345e+17, 1.288744324452407e+17, 1.288744324493033e+17, 1.288744324532095e+17, 1.288744324572719e+17, 1.288744324613345e+17, 1.288744324652407e+17, 1.288744324693033e+17, 1.288744324732095e+17, 1.288744324772721e+17, 1.288744324813345e+17, 1.288744324852408e+17, 1.288744324893033e+17, 1.288744324932095e+17, 1.288744324972721e+17, 1.288744325013344e+17, 1.288744325052407e+17, 1.288744325093033e+17, 1.288744325132095e+17, 1.288744325172721e+17, 1.288744325213345e+17, 1.288744325252408e+17, 1.288744325293032e+17, 1.288744325332095e+17, 1.288744325372721e+17, 1.288744325413344e+17, 1.288744325452408e+17, 1.288744325493032e+17, 1.288744325532095e+17, 1.288744325572719e+17, 1.288744325613345e+17, 1.288744325652408e+17, 1.288744325693032e+17, 1.288744325732096e+17, 1.288744325772719e+17, 1.288744325813345e+17, 1.288744325852407e+17, 1.288744325893032e+17, 1.288744325932095e+17, 1.288744325972719e+17, 1.288744326013345e+17, 1.288744326052407e+17, 1.288744326093033e+17, 1.288744326132095e+17, 1.288744326172719e+17, 1.288744326213345e+17, 1.288744326252407e+17, 1.288744326293032e+17, 1.288744326332095e+17, 1.288744326372719e+17, 1.288744326413345e+17, 1.288744326452407e+17, 1.288744326493033e+17, 1.288744326532095e+17, 1.288744326572721e+17, 1.288744326613345e+17, 1.288744326652407e+17, 1.288744326693033e+17, 1.288744326732095e+17, 1.288744326772719e+17, 1.288744326813345e+17, 1.288744326852407e+17, 1.288744326893033e+17, 1.288744326932095e+17, 1.288744326972721e+17, 1.288744327013345e+17, 1.288744327052407e+17, 1.288744327093033e+17, 1.288744327132095e+17, 1.288744327172721e+17, 1.288744327213345e+17, 1.288744327252407e+17, 1.288744327293033e+17, 1.288744327332095e+17, 1.288744327372721e+17, 1.288744327413345e+17, 1.288744327452408e+17, 1.288744327493033e+17, 1.288744327532095e+17, 1.288744327572721e+17, 1.288744327613344e+17, 1.288744327652407e+17, 1.288744327693033e+17, 1.288744327732095e+17, 1.288744327772721e+17, 1.288744327813345e+17, 1.288744327852408e+17, 1.288744327893032e+17, 1.288744327932095e+17, 1.288744327972721e+17, 1.288744328013344e+17, 1.288744328052408e+17, 1.288744328093032e+17, 1.288744328132095e+17, 1.288744328172719e+17, 1.288744328213345e+17, 1.288744328252408e+17, 1.288744328293032e+17, 1.288744328332096e+17, 1.288744328372719e+17, 1.288744328413345e+17, 1.288744328452407e+17, 1.288744328493032e+17, 1.288744328532095e+17, 1.288744328572719e+17, 1.288744328613345e+17, 1.288744328652407e+17, 1.288744328693033e+17, 1.288744328732095e+17, 1.288744328772719e+17, 1.288744328813345e+17, 1.288744328852407e+17, 1.288744328893032e+17, 1.288744328932095e+17, 1.288744328972719e+17, 1.288744329013345e+17, 1.288744329052407e+17, 1.288744329093033e+17, 1.288744329132095e+17, 1.288744329172721e+17, 1.288744329213345e+17, 1.288744329252407e+17, 1.288744329293033e+17, 1.288744329332095e+17, 1.288744329372719e+17, 1.288744329413345e+17, 1.288744329452407e+17, 1.288744329493033e+17, 1.288744329532095e+17, 1.288744329572721e+17, 1.288744329613345e+17, 1.288744329652407e+17, 1.288744329693033e+17, 1.288744329732095e+17, 1.288744329772721e+17, 1.288744329813345e+17, 1.288744329852407e+17, 1.288744329893033e+17, 1.288744329932095e+17, 1.288744329972721e+17, 1.288744330013344e+17, 1.288744330052408e+17, 1.288744330093033e+17, 1.288744330132095e+17, 1.288744330172721e+17, 1.288744330213344e+17, 1.288744330252407e+17, 1.288744330293032e+17, 1.288744330332095e+17, 1.288744330372721e+17, 1.288744330413345e+17, 1.288744330452408e+17, 1.288744330493032e+17, 1.288744330532096e+17, 1.288744330572719e+17, 1.288744330613344e+17, 1.288744330652408e+17, 1.288744330693032e+17, 1.288744330732095e+17, 1.288744330772719e+17, 1.288744330813345e+17, 1.288744330852407e+17, 1.288744330893033e+17, 1.288744330932096e+17, 1.288744330972719e+17, 1.288744331013345e+17, 1.288744331052407e+17, 1.288744331093032e+17, 1.288744331132095e+17, 1.288744331172719e+17, 1.288744331213345e+17, 1.288744331252407e+17, 1.288744331293033e+17, 1.288744331332095e+17, 1.288744331372719e+17, 1.288744331413345e+17, 1.288744331452407e+17, 1.288744331493032e+17, 1.288744331532095e+17, 1.288744331572719e+17, 1.288744331613345e+17, 1.288744331652407e+17, 1.288744331693033e+17, 1.288744331732095e+17, 1.288744331772721e+17, 1.288744331813345e+17, 1.288744331852407e+17, 1.288744331893033e+17, 1.288744331932095e+17, 1.288744331972719e+17, 1.288744332013345e+17, 1.288744332052407e+17, 1.288744332093033e+17, 1.288744332132095e+17, 1.288744332172721e+17, 1.288744332213345e+17, 1.288744332252407e+17, 1.288744332293033e+17, 1.288744332332095e+17, 1.288744332372721e+17, 1.288744332413345e+17, 1.288744332452407e+17, 1.288744332493033e+17, 1.288744332532095e+17, 1.288744332572721e+17, 1.288744332613344e+17, 1.288744332652408e+17, 1.288744332693033e+17, 1.288744332732095e+17, 1.288744332772721e+17, 1.288744332813344e+17, 1.288744332852407e+17, 1.288744332893032e+17, 1.288744332932095e+17, 1.288744332972721e+17, 1.288744333013345e+17, 1.288744333052408e+17, 1.288744333093032e+17, 1.288744333132096e+17, 1.288744333172719e+17, 1.288744333213344e+17, 1.288744333252408e+17, 1.288744333293032e+17, 1.288744333332095e+17, 1.288744333372719e+17, 1.288744333413345e+17, 1.288744333452407e+17, 1.288744333493033e+17, 1.288744333532096e+17, 1.288744333572719e+17, 1.288744333613345e+17, 1.288744333652407e+17, 1.288744333693032e+17, 1.288744333732095e+17, 1.288744333772719e+17, 1.288744333813345e+17, 1.288744333852407e+17, 1.288744333893033e+17, 1.288744333932095e+17, 1.288744333972719e+17, 1.288744334013345e+17, 1.288744334052407e+17, 1.288744334093033e+17, 1.288744334132095e+17, 1.288744334172719e+17, 1.288744334213345e+17, 1.288744334252407e+17, 1.288744334293033e+17, 1.288744334332095e+17, 1.288744334372721e+17, 1.288744334413345e+17, 1.288744334452407e+17, 1.288744334493033e+17, 1.288744334532095e+17, 1.288744334572719e+17, 1.288744334613345e+17, 1.288744334652407e+17, 1.288744334693033e+17, 1.288744334732095e+17, 1.288744334772721e+17, 1.288744334813345e+17, 1.288744334852407e+17, 1.288744334893033e+17, 1.288744334932095e+17, 1.288744334972721e+17, 1.288744335013345e+17, 1.288744335052407e+17, 1.288744335093033e+17, 1.288744335132095e+17, 1.288744335172721e+17, 1.288744335213344e+17, 1.288744335252408e+17, 1.288744335293033e+17, 1.288744335332095e+17, 1.288744335372721e+17, 1.288744335413344e+17, 1.288744335452407e+17, 1.288744335493032e+17, 1.288744335532095e+17, 1.288744335572721e+17, 1.288744335613345e+17, 1.288744335652408e+17, 1.288744335693032e+17, 1.288744335732096e+17, 1.288744335772719e+17, 1.288744335813344e+17, 1.288744335852408e+17, 1.288744335893032e+17, 1.288744335932095e+17, 1.288744335972719e+17, 1.288744336013345e+17, 1.288744336052407e+17, 1.288744336093033e+17, 1.288744336132096e+17, 1.288744336172719e+17, 1.288744336213345e+17, 1.288744336252407e+17, 1.288744336293032e+17, 1.288744336332095e+17, 1.288744336372719e+17, 1.288744336413345e+17, 1.288744336452407e+17, 1.288744336493033e+17, 1.288744336532095e+17, 1.288744336572719e+17, 1.288744336613345e+17, 1.288744336652407e+17, 1.288744336693033e+17, 1.288744336732095e+17, 1.288744336772719e+17, 1.288744336813345e+17, 1.288744336852407e+17, 1.288744336893033e+17, 1.288744336932095e+17, 1.288744336972721e+17, 1.288744337013345e+17, 1.288744337052407e+17, 1.288744337093033e+17, 1.288744337132095e+17, 1.288744337172719e+17, 1.288744337213345e+17, 1.288744337252407e+17, 1.288744337293033e+17, 1.288744337332095e+17, 1.288744337372721e+17, 1.288744337413345e+17, 1.288744337452408e+17, 1.288744337493033e+17, 1.288744337532095e+17, 1.288744337572721e+17, 1.288744337613344e+17, 1.288744337652407e+17, 1.288744337706632e+17, 1.288744337745696e+17, 1.288744337786319e+17, 1.288744337826944e+17, 1.288744337866008e+17, 1.288744337906632e+17, 1.288744337945696e+17, 1.288744337986319e+17, 1.288744338026945e+17, 1.288744338066007e+17, 1.288744338106632e+17, 1.288744338145696e+17, 1.288744338186319e+17, 1.288744338226945e+17, 1.288744338266007e+17, 1.288744338306632e+17, 1.288744338345695e+17, 1.288744338386319e+17, 1.288744338426945e+17, 1.288744338466007e+17, 1.288744338506633e+17, 1.288744338545695e+17, 1.288744338586319e+17, 1.288744338626945e+17, 1.288744338666007e+17, 1.288744338706632e+17, 1.288744338745695e+17, 1.288744338786319e+17, 1.288744338826945e+17, 1.288744338866007e+17, 1.288744338906633e+17, 1.288744338945695e+17, 1.288744338986321e+17, 1.288744339026945e+17, 1.288744339066007e+17, 1.288744339106633e+17, 1.288744339145695e+17, 1.288744339186319e+17, 1.288744339226945e+17, 1.288744339266007e+17, 1.288744339306633e+17, 1.288744339345695e+17, 1.288744339386321e+17, 1.288744339426945e+17, 1.288744339466008e+17, 1.288744339506633e+17, 1.288744339545695e+17, 1.288744339586321e+17, 1.288744339626945e+17, 1.288744339666007e+17, 1.288744339706633e+17, 1.288744339745695e+17, 1.288744339786321e+17, 1.288744339826944e+17, 1.288744339866008e+17, 1.288744339906633e+17, 1.288744339945696e+17, 1.288744339986321e+17, 1.288744340026944e+17, 1.288744340066008e+17, 1.288744340106632e+17, 1.288744340145695e+17, 1.288744340186321e+17, 1.288744340226945e+17, 1.288744340266008e+17, 1.288744340306632e+17, 1.288744340345696e+17, 1.288744340386319e+17, 1.288744340426944e+17, 1.288744340466008e+17, 1.288744340506632e+17, 1.288744340545696e+17, 1.288744340586319e+17, 1.288744340626945e+17, 1.288744340666007e+17, 1.288744340706633e+17, 1.288744340745696e+17, 1.288744340786319e+17, 1.288744340826945e+17, 1.288744340866007e+17, 1.288744340906632e+17, 1.288744340945695e+17, 1.288744340986319e+17, 1.288744341026945e+17, 1.288744341066007e+17, 1.288744341106633e+17, 1.288744341145695e+17, 1.288744341186319e+17, 1.288744341226945e+17, 1.288744341266007e+17, 1.288744341306633e+17, 1.288744341345695e+17, 1.288744341386319e+17, 1.288744341426945e+17, 1.288744341466007e+17, 1.288744341506633e+17, 1.288744341545695e+17, 1.288744341586321e+17, 1.288744341626945e+17, 1.288744341666008e+17, 1.288744341706633e+17, 1.288744341745695e+17, 1.288744341786319e+17, 1.288744341826945e+17, 1.288744341866007e+17, 1.288744341906633e+17, 1.288744341945695e+17, 1.288744341986321e+17, 1.288744342026945e+17, 1.288744342066008e+17, 1.288744342106633e+17, 1.288744342145695e+17, 1.288744342186321e+17, 1.288744342226945e+17, 1.288744342266007e+17, 1.288744342306633e+17, 1.288744342345695e+17, 1.288744342386321e+17, 1.288744342426944e+17, 1.288744342466008e+17, 1.288744342506633e+17, 1.288744342545696e+17, 1.288744342586321e+17, 1.288744342626944e+17, 1.288744342666008e+17, 1.288744342706632e+17, 1.288744342745695e+17, 1.288744342786321e+17, 1.288744342826945e+17, 1.288744342866008e+17, 1.288744342906632e+17, 1.288744342945696e+17, 1.288744342986319e+17, 1.288744343026944e+17, 1.288744343066008e+17, 1.288744343106632e+17, 1.288744343145696e+17, 1.288744343186319e+17, 1.288744343226945e+17, 1.288744343266007e+17, 1.288744343306633e+17, 1.288744343345696e+17, 1.288744343386319e+17, 1.288744343426945e+17, 1.288744343466007e+17, 1.288744343506632e+17, 1.288744343545695e+17, 1.288744343586319e+17, 1.288744343626945e+17, 1.288744343666007e+17, 1.288744343706633e+17, 1.288744343745695e+17, 1.288744343786319e+17, 1.288744343826945e+17, 1.288744343866007e+17, 1.288744343906633e+17, 1.288744343945695e+17, 1.288744343986319e+17, 1.288744344026945e+17, 1.288744344066007e+17, 1.288744344106633e+17, 1.288744344145695e+17, 1.288744344186321e+17, 1.288744344226945e+17, 1.288744344266008e+17, 1.288744344306633e+17, 1.288744344345695e+17, 1.288744344386319e+17, 1.288744344426945e+17, 1.288744344466007e+17, 1.288744344506633e+17, 1.288744344545695e+17, 1.288744344586321e+17, 1.288744344626945e+17, 1.288744344666008e+17, 1.288744344706633e+17, 1.288744344745695e+17, 1.288744344786321e+17, 1.288744344826944e+17, 1.288744344866008e+17, 1.288744344906633e+17, 1.288744344945695e+17, 1.288744344986321e+17, 1.288744345026945e+17, 1.288744345066008e+17, 1.288744345106632e+17, 1.288744345145696e+17, 1.288744345186321e+17, 1.288744345226944e+17, 1.288744345266008e+17, 1.288744345306632e+17, 1.288744345345695e+17, 1.288744345386319e+17, 1.288744345426945e+17, 1.288744345466008e+17, 1.288744345506632e+17, 1.288744345545696e+17, 1.288744345586319e+17, 1.288744345626944e+17, 1.288744345666007e+17, 1.288744345706632e+17, 1.288744345745696e+17, 1.288744345786319e+17, 1.288744345826945e+17, 1.288744345866007e+17, 1.288744345906633e+17, 1.288744345945695e+17, 1.288744345986319e+17, 1.288744346026945e+17, 1.288744346066007e+17, 1.288744346106632e+17, 1.288744346145695e+17, 1.288744346186319e+17, 1.288744346226945e+17, 1.288744346266007e+17, 1.288744346306633e+17, 1.288744346345695e+17, 1.288744346386319e+17, 1.288744346426945e+17, 1.288744346466007e+17, 1.288744346506633e+17, 1.288744346545695e+17, 1.288744346586319e+17, 1.288744346626945e+17, 1.288744346666007e+17, 1.288744346706633e+17, 1.288744346745695e+17, 1.288744346786321e+17, 1.288744346826945e+17, 1.288744346866008e+17, 1.288744346906633e+17, 1.288744346945695e+17, 1.288744346986319e+17, 1.288744347026945e+17, 1.288744347066007e+17, 1.288744347106633e+17, 1.288744347145695e+17, 1.288744347186321e+17, 1.288744347226945e+17, 1.288744347266008e+17, 1.288744347306633e+17, 1.288744347345695e+17, 1.288744347386321e+17, 1.288744347426944e+17, 1.288744347466008e+17, 1.288744347506633e+17, 1.288744347545695e+17, 1.288744347586321e+17, 1.288744347626945e+17, 1.288744347666008e+17, 1.288744347706632e+17, 1.288744347745696e+17, 1.288744347786321e+17, 1.288744347826944e+17, 1.288744347866008e+17, 1.288744347906632e+17, 1.288744347945695e+17, 1.288744347986319e+17, 1.288744348026945e+17, 1.288744348066008e+17, 1.288744348106632e+17, 1.288744348145696e+17, 1.288744348186319e+17, 1.288744348226945e+17, 1.288744348266007e+17, 1.288744348306632e+17, 1.288744348345696e+17, 1.288744348386319e+17, 1.288744348426945e+17, 1.288744348466007e+17, 1.288744348506633e+17, 1.288744348545695e+17, 1.288744348586319e+17, 1.288744348626945e+17, 1.288744348666007e+17, 1.288744348706632e+17, 1.288744348745695e+17, 1.288744348786319e+17, 1.288744348826945e+17, 1.288744348866007e+17, 1.288744348906633e+17, 1.288744348945695e+17, 1.288744348986319e+17, 1.288744349026945e+17, 1.288744349066007e+17, 1.288744349106633e+17, 1.288744349145695e+17, 1.288744349186319e+17, 1.288744349226945e+17, 1.288744349266007e+17, 1.288744349306633e+17, 1.288744349345695e+17, 1.288744349386321e+17, 1.288744349426945e+17, 1.288744349466008e+17, 1.288744349506633e+17, 1.288744349545695e+17, 1.288744349586319e+17, 1.288744349626945e+17, 1.288744349666007e+17, 1.288744349706633e+17, 1.288744349745695e+17, 1.288744349786321e+17, 1.288744349826945e+17, 1.288744349866008e+17, 1.288744349906633e+17, 1.288744349945695e+17, 1.288744349986321e+17, 1.288744350026944e+17, 1.288744350066008e+17, 1.288744350106633e+17, 1.288744350145695e+17, 1.288744350186321e+17, 1.288744350226945e+17, 1.288744350266008e+17, 1.288744350306632e+17, 1.288744350345696e+17},
			             {1.288743885967732e+17, 1.288743886008357e+17, 1.288743886048983e+17, 1.288743886088045e+17, 1.288743886128671e+17, 1.288743886167732e+17, 1.288743886208358e+17},
			             {1.288744002332096e+17, 1.288744002372719e+17, 1.288744002413345e+17, 1.288744002452407e+17, 1.288744002493032e+17, 1.288744002532095e+17, 1.288744002572719e+17, 1.288744002613345e+17, 1.288744002652407e+17, 1.288744002693033e+17, 1.288744002732095e+17, 1.288744002772719e+17, 1.288744002813345e+17, 1.288744002852407e+17, 1.288744002893032e+17, 1.288744002932095e+17, 1.288744002972719e+17, 1.288744003013345e+17, 1.288744003052407e+17, 1.288744003093033e+17, 1.288744003132095e+17, 1.288744003172721e+17, 1.288744003213345e+17, 1.288744003252407e+17, 1.288744003293033e+17, 1.288744003332095e+17, 1.288744003372719e+17, 1.288744003413345e+17, 1.288744003452407e+17, 1.288744003532095e+17, 1.288744003572721e+17, 1.288744003613345e+17, 1.288744003652407e+17, 1.288744003693033e+17, 1.288744003732095e+17, 1.288744003772721e+17, 1.288744003813345e+17, 1.288744003852407e+17, 1.288744003893033e+17, 1.288744003932095e+17, 1.288744003972721e+17, 1.288744004013344e+17, 1.288744004052408e+17, 1.288744004093033e+17, 1.288744004132095e+17, 1.288744004172721e+17, 1.288744004213344e+17, 1.288744004252407e+17, 1.288744004293032e+17, 1.288744004332095e+17, 1.288744004452408e+17, 1.288744004532096e+17, 1.288744004572719e+17, 1.288744004613344e+17, 1.288744004652408e+17},
			             {1.288744007613345e+17, 1.288744007652407e+17, 1.288744007693032e+17, 1.288744007732095e+17, 1.288744007772719e+17, 1.288744007813345e+17, 1.288744007852407e+17, 1.288744007893033e+17, 1.288744007932095e+17, 1.288744007972719e+17, 1.288744008013345e+17, 1.288744008052407e+17, 1.288744008093033e+17, 1.288744008132095e+17, 1.288744008172719e+17, 1.288744008213345e+17, 1.288744008252407e+17, 1.288744008293033e+17, 1.288744008332095e+17, 1.288744008372721e+17, 1.288744008413345e+17, 1.288744008452407e+17, 1.288744008493033e+17, 1.288744008532095e+17, 1.288744008572719e+17, 1.288744008613345e+17, 1.288744008652407e+17, 1.288744008693033e+17, 1.288744008732095e+17, 1.288744008772721e+17, 1.288744008813345e+17, 1.288744008852408e+17, 1.288744008893033e+17, 1.288744008932095e+17, 1.288744008972721e+17, 1.288744009013345e+17, 1.288744009052407e+17, 1.288744009093033e+17, 1.288744009132095e+17, 1.288744009172721e+17, 1.288744009213345e+17, 1.288744009252408e+17, 1.288744009293033e+17, 1.288744009332095e+17, 1.288744009372721e+17, 1.288744009413344e+17, 1.288744009452407e+17, 1.288744009493032e+17, 1.288744009532095e+17, 1.288744009572721e+17, 1.288744009613345e+17, 1.288744009652408e+17, 1.288744009693032e+17, 1.288744009732096e+17, 1.288744009772719e+17, 1.288744009813344e+17, 1.288744009852408e+17, 1.288744009893032e+17, 1.288744009932095e+17, 1.288744009972719e+17, 1.288744010013345e+17, 1.288744010052407e+17, 1.288744010093033e+17, 1.288744010132096e+17, 1.288744010172719e+17, 1.288744010213345e+17, 1.288744010252407e+17, 1.288744010293032e+17, 1.288744010332095e+17, 1.288744010372719e+17, 1.288744010413345e+17, 1.288744010452407e+17},
			             {1.288743983413345e+17, 1.288743983452407e+17, 1.288743983493033e+17, 1.288743983532095e+17, 1.288743983572721e+17, 1.288743983613344e+17, 1.288743983652408e+17},
			             {1.288744015493032e+17, 1.288744015532095e+17, 1.288744015572719e+17, 1.288744015613345e+17, 1.288744015652407e+17, 1.288744015693033e+17, 1.288744015732095e+17},
			             {1.288744027893033e+17, 1.288744027932096e+17, 1.288744027972719e+17, 1.288744028013345e+17, 1.288744028052407e+17},
			             {1.288744028013345e+17, 1.288744028052407e+17, 1.288744028093032e+17, 1.288744028132095e+17, 1.288744028172719e+17, 1.288744028213345e+17, 1.288744028252407e+17, 1.288744028293033e+17},
			             {1.288743950888045e+17, 1.288743950928669e+17, 1.288743950967732e+17, 1.288743951008357e+17, 1.288743951048983e+17, 1.288743951088045e+17, 1.288743951128669e+17},
			             {1.288743916728671e+17, 1.288743916767732e+17, 1.288743916808357e+17, 1.288743916848982e+17, 1.288743916888045e+17, 1.288743916928671e+17, 1.288743916967732e+17},
			             {1.288743920767732e+17, 1.288743920808357e+17, 1.288743920848983e+17, 1.288743920888045e+17, 1.288743920928671e+17},
			             {1.288743937888046e+17, 1.288743937928669e+17, 1.288743937967732e+17, 1.288743938008357e+17, 1.288743938048982e+17, 1.288743938088045e+17},
			             {1.288743978813345e+17, 1.288743978852408e+17, 1.288743978893032e+17, 1.288743978932095e+17, 1.288743978972721e+17, 1.288743979013344e+17},
			             {1.288743952208358e+17, 1.288743952248983e+17, 1.288743952288045e+17, 1.288743952328671e+17, 1.288743952367732e+17},
			             {1.288744063852407e+17, 1.288744063893033e+17, 1.288744063932095e+17, 1.288744063972719e+17, 1.288744064013345e+17, 1.288744064052407e+17, 1.288744064093033e+17, 1.288744064132095e+17, 1.288744064172719e+17, 1.288744064213345e+17, 1.288744064252407e+17, 1.288744064293033e+17, 1.288744064332095e+17, 1.288744064372721e+17, 1.288744064413345e+17, 1.288744064452407e+17, 1.288744064493033e+17},
			             {1.288744086532096e+17, 1.288744086572719e+17, 1.288744086613345e+17, 1.288744086652407e+17, 1.288744086693032e+17, 1.288744086732095e+17, 1.288744086772719e+17, 1.288744086813345e+17, 1.288744086852407e+17, 1.288744086893033e+17, 1.288744086932095e+17, 1.288744086972719e+17, 1.288744087013345e+17, 1.288744087052407e+17, 1.288744087093033e+17, 1.288744087132095e+17, 1.288744087172719e+17, 1.288744087213345e+17, 1.288744087252407e+17, 1.288744087293033e+17, 1.288744087332095e+17, 1.288744087372721e+17, 1.288744087413345e+17},
			             {1.288744090372721e+17, 1.288744090413345e+17, 1.288744090452408e+17, 1.288744090493033e+17, 1.288744090532095e+17, 1.288744090572721e+17, 1.288744090613344e+17, 1.288744090652407e+17, 1.288744090693033e+17, 1.288744090732095e+17, 1.288744090772721e+17, 1.288744090813345e+17, 1.288744090852408e+17, 1.288744090893032e+17, 1.288744090932095e+17, 1.288744090972721e+17, 1.288744091013344e+17, 1.288744091052408e+17, 1.288744091093032e+17, 1.288744091132095e+17, 1.288744091172719e+17, 1.288744091213345e+17, 1.288744091252408e+17, 1.288744091293032e+17, 1.288744091332096e+17, 1.288744091372719e+17, 1.288744091413345e+17, 1.288744091452407e+17, 1.288744091493032e+17, 1.288744091532095e+17, 1.288744091572719e+17, 1.288744091613345e+17, 1.288744091652407e+17, 1.288744091693033e+17, 1.288744091732095e+17, 1.288744091772719e+17, 1.288744091813345e+17, 1.288744091852407e+17, 1.288744091893032e+17, 1.288744091932095e+17, 1.288744091972719e+17, 1.288744092013345e+17, 1.288744092052407e+17, 1.288744092093033e+17, 1.288744092132095e+17, 1.288744092172721e+17, 1.288744092213345e+17},
			             {1.288744092893033e+17, 1.288744092932095e+17, 1.288744092972721e+17, 1.288744093013345e+17, 1.288744093052408e+17, 1.288744093093033e+17, 1.288744093132095e+17, 1.288744093172721e+17, 1.288744093213344e+17, 1.288744093252407e+17, 1.288744093293033e+17, 1.288744093332095e+17, 1.288744093372721e+17, 1.288744093413345e+17, 1.288744093452408e+17, 1.288744093493032e+17, 1.288744093532095e+17},
			             {1.288744094052407e+17, 1.288744094093032e+17, 1.288744094132095e+17, 1.288744094172719e+17, 1.288744094213345e+17, 1.288744094252407e+17, 1.288744094293033e+17, 1.288744094332095e+17, 1.288744094372719e+17, 1.288744094413345e+17, 1.288744094452407e+17, 1.288744094493032e+17},
			             {1.288744097732095e+17, 1.288744097772721e+17, 1.288744097813345e+17, 1.288744097852407e+17, 1.288744097893033e+17, 1.288744097932095e+17, 1.288744097972721e+17, 1.288744098013345e+17, 1.288744098052407e+17, 1.288744098093033e+17, 1.288744098132095e+17, 1.288744098172721e+17, 1.288744098213344e+17, 1.288744098252408e+17, 1.288744098293033e+17, 1.288744098332095e+17},
			             {1.288744098372721e+17, 1.288744098413344e+17, 1.288744098452407e+17, 1.288744098493032e+17, 1.288744098532095e+17},
			             {1.288744108413344e+17, 1.288744108452407e+17, 1.288744108493033e+17, 1.288744108532095e+17, 1.288744108572721e+17, 1.288744108613345e+17},
			             {1.288744109572719e+17, 1.288744109613345e+17, 1.288744109652407e+17, 1.288744109693032e+17, 1.288744109732095e+17, 1.288744109772719e+17, 1.288744109813345e+17, 1.288744109852407e+17, 1.288744109893033e+17},
			             {1.288744121532095e+17, 1.288744121572721e+17, 1.288744121613345e+17, 1.288744121652408e+17, 1.288744121693032e+17, 1.288744121732096e+17, 1.288744121772719e+17, 1.288744121813344e+17, 1.288744121852408e+17, 1.288744121893032e+17, 1.288744121932095e+17, 1.288744121972719e+17, 1.288744122013345e+17, 1.288744122052407e+17, 1.288744122093033e+17, 1.288744122132096e+17, 1.288744122172719e+17, 1.288744122213345e+17, 1.288744122252407e+17, 1.288744122293032e+17, 1.288744122332095e+17, 1.288744122372719e+17, 1.288744122413345e+17, 1.288744122452407e+17, 1.288744122493033e+17, 1.288744122532095e+17, 1.288744122572719e+17, 1.288744122613345e+17},
			             {1.288744126052408e+17, 1.288744126093033e+17, 1.288744126132095e+17, 1.288744126172721e+17, 1.288744126213344e+17, 1.288744126252407e+17, 1.288744126293033e+17, 1.288744126332095e+17, 1.288744126372721e+17, 1.288744126413345e+17, 1.288744126452408e+17, 1.288744126493032e+17, 1.288744126532095e+17, 1.288744126572721e+17, 1.288744126613344e+17, 1.288744126652408e+17},
			             {1.288744146132095e+17, 1.288744146172719e+17, 1.288744146213345e+17, 1.288744146252407e+17, 1.288744146293033e+17, 1.288744146332095e+17, 1.288744146372721e+17, 1.288744146413345e+17, 1.288744146452408e+17, 1.288744146493033e+17, 1.288744146532095e+17, 1.288744146572721e+17, 1.288744146613344e+17},
			             {1.288744155013345e+17, 1.288744155052408e+17, 1.288744155093032e+17, 1.288744155132096e+17, 1.288744155172719e+17, 1.288744155213345e+17, 1.288744155252407e+17, 1.288744155293032e+17, 1.288744155332095e+17, 1.288744155372719e+17, 1.288744155413345e+17, 1.288744155452407e+17, 1.288744155493033e+17, 1.288744155532095e+17, 1.288744155572719e+17, 1.288744155613345e+17, 1.288744155652407e+17, 1.288744155693032e+17, 1.288744155732095e+17, 1.288744155772719e+17, 1.288744155813345e+17, 1.288744155852407e+17},
			             {1.288744167013344e+17, 1.288744167052407e+17, 1.288744167093033e+17, 1.288744167132095e+17, 1.288744167172721e+17, 1.288744167213345e+17, 1.288744167252408e+17, 1.288744167293032e+17, 1.288744167332095e+17},
			             {1.288744176413345e+17, 1.288744176452407e+17, 1.288744176493033e+17, 1.288744176532095e+17, 1.288744176572719e+17, 1.288744176613345e+17, 1.288744176652407e+17, 1.288744176693033e+17, 1.288744176732095e+17, 1.288744176772721e+17, 1.288744176813345e+17, 1.288744176852407e+17, 1.288744176893033e+17, 1.288744176932095e+17},
			             {1.288744204693033e+17, 1.288744204732095e+17, 1.288744204772719e+17, 1.288744204813345e+17, 1.288744204852407e+17, 1.288744204893033e+17, 1.288744204932095e+17, 1.288744204972721e+17, 1.288744205013345e+17, 1.288744205052408e+17, 1.288744205093033e+17, 1.288744205132095e+17, 1.288744205172721e+17, 1.288744205213344e+17},
			             {1.288744161693033e+17, 1.288744161732095e+17, 1.288744161772721e+17, 1.288744161813345e+17, 1.288744161852407e+17, 1.288744161893033e+17, 1.288744161932095e+17, 1.288744161972721e+17},
			             {1.288744217893033e+17, 1.288744217932095e+17, 1.288744217972721e+17, 1.288744218013344e+17, 1.288744218052408e+17, 1.288744218093033e+17, 1.288744218132095e+17, 1.288744218172721e+17, 1.288744218213344e+17, 1.288744218252407e+17, 1.288744218293032e+17, 1.288744218332095e+17},
			             {1.288744282172719e+17, 1.288744282213345e+17, 1.288744282252408e+17, 1.288744282293032e+17, 1.288744282332096e+17, 1.288744282372719e+17, 1.288744282413345e+17, 1.288744282452407e+17, 1.288744282493032e+17, 1.288744282532095e+17},
			             {1.288744225452408e+17, 1.288744225493033e+17, 1.288744225532095e+17, 1.288744225572721e+17, 1.288744225613344e+17, 1.288744225652407e+17, 1.288744225693033e+17, 1.288744225732095e+17, 1.288744225772721e+17, 1.288744225813345e+17},
			             {1.288744270813345e+17, 1.288744270852407e+17, 1.288744270893033e+17, 1.288744270932095e+17, 1.288744270972721e+17, 1.288744271013345e+17, 1.288744271052407e+17, 1.288744271093033e+17, 1.288744271132095e+17, 1.288744271172721e+17},
			             {1.288744305213345e+17, 1.288744305252408e+17, 1.288744305293032e+17, 1.288744305332096e+17, 1.288744305372719e+17, 1.288744305413345e+17, 1.288744305452407e+17, 1.288744305493032e+17},
			             {1.288744255413345e+17, 1.288744255452407e+17, 1.288744255493033e+17, 1.288744255532095e+17, 1.288744255572719e+17, 1.288744255613345e+17, 1.288744255652407e+17, 1.288744255693033e+17, 1.288744255732095e+17, 1.288744255772721e+17, 1.288744255813345e+17, 1.288744255852407e+17, 1.288744255893033e+17, 1.288744255932095e+17, 1.288744255972721e+17, 1.288744256013345e+17, 1.288744256052407e+17, 1.288744256093033e+17, 1.288744256132095e+17, 1.288744256172721e+17, 1.288744256213344e+17, 1.288744256252408e+17, 1.288744256293033e+17, 1.288744256332095e+17, 1.288744256372721e+17, 1.288744256413344e+17, 1.288744256452407e+17, 1.288744256493032e+17, 1.288744256532095e+17, 1.288744256572721e+17, 1.288744256613345e+17, 1.288744256652408e+17, 1.288744256693032e+17, 1.288744256732096e+17, 1.288744256772719e+17},
			             {1.288744256932095e+17, 1.288744256972719e+17, 1.288744257013345e+17, 1.288744257052407e+17, 1.288744257093033e+17, 1.288744257132096e+17, 1.288744257172719e+17, 1.288744257213345e+17, 1.288744257252407e+17, 1.288744257293032e+17, 1.288744257332095e+17, 1.288744257372719e+17, 1.288744257413345e+17, 1.288744257452407e+17, 1.288744257493033e+17, 1.288744257532095e+17, 1.288744257572719e+17, 1.288744257613345e+17, 1.288744257652407e+17, 1.288744257693033e+17, 1.288744257732095e+17, 1.288744257772719e+17, 1.288744257813345e+17, 1.288744257852407e+17, 1.288744257893033e+17, 1.288744257932095e+17, 1.288744257972721e+17, 1.288744258013345e+17, 1.288744258052407e+17, 1.288744258093033e+17, 1.288744258132095e+17, 1.288744258172719e+17, 1.288744258213345e+17, 1.288744258252407e+17, 1.288744258293033e+17, 1.288744258332095e+17, 1.288744258372721e+17, 1.288744258413345e+17, 1.288744258452407e+17, 1.288744258493033e+17, 1.288744258532095e+17, 1.288744258572721e+17, 1.288744258613345e+17, 1.288744258652407e+17, 1.288744258693033e+17, 1.288744258732095e+17, 1.288744258772721e+17, 1.288744258813345e+17, 1.288744258852408e+17, 1.288744258893033e+17, 1.288744258932095e+17, 1.288744258972721e+17, 1.288744259013344e+17, 1.288744259052407e+17, 1.288744259093032e+17, 1.288744259132095e+17, 1.288744259172721e+17, 1.288744259213345e+17, 1.288744259252408e+17, 1.288744259293032e+17, 1.288744259332096e+17, 1.288744259372719e+17, 1.288744259413344e+17, 1.288744259452408e+17, 1.288744259493032e+17, 1.288744259532095e+17, 1.288744259572719e+17, 1.288744259613345e+17, 1.288744259652407e+17, 1.288744259693033e+17, 1.288744259732096e+17, 1.288744259772719e+17, 1.288744259813345e+17, 1.288744259852407e+17, 1.288744259893032e+17, 1.288744259932095e+17, 1.288744259972719e+17, 1.288744260013345e+17, 1.288744260052407e+17, 1.288744260093033e+17, 1.288744260132095e+17, 1.288744260172719e+17, 1.288744260213345e+17, 1.288744260252407e+17, 1.288744260293033e+17, 1.288744260332095e+17, 1.288744260372719e+17, 1.288744260413345e+17, 1.288744260452407e+17, 1.288744260493033e+17, 1.288744260532095e+17, 1.288744260572721e+17, 1.288744260613345e+17, 1.288744260652407e+17, 1.288744260693033e+17, 1.288744260732095e+17, 1.288744260772719e+17, 1.288744260813345e+17, 1.288744260852407e+17, 1.288744260893033e+17, 1.288744260932095e+17, 1.288744260972721e+17, 1.288744261013345e+17, 1.288744261052408e+17, 1.288744261093033e+17, 1.288744261132095e+17, 1.288744261172721e+17, 1.288744261213344e+17, 1.288744261252407e+17, 1.288744261293033e+17, 1.288744261332095e+17, 1.288744261372721e+17, 1.288744261413345e+17, 1.288744261452408e+17, 1.288744261493032e+17, 1.288744261532095e+17, 1.288744261572721e+17, 1.288744261613344e+17, 1.288744261652408e+17, 1.288744261693032e+17, 1.288744261732095e+17, 1.288744261772719e+17, 1.288744261813345e+17, 1.288744261852408e+17, 1.288744261893032e+17, 1.288744261932096e+17, 1.288744261972719e+17, 1.288744262013345e+17, 1.288744262052407e+17, 1.288744262093032e+17, 1.288744262132095e+17, 1.288744262172719e+17, 1.288744262213345e+17, 1.288744262252407e+17, 1.288744262293033e+17, 1.288744262332095e+17, 1.288744262372719e+17, 1.288744262413345e+17, 1.288744262452407e+17, 1.288744262493032e+17, 1.288744262532095e+17, 1.288744262572719e+17, 1.288744262613345e+17, 1.288744262652407e+17, 1.288744262693033e+17, 1.288744262732095e+17, 1.288744262772719e+17, 1.288744262813345e+17, 1.288744262852407e+17, 1.288744262893033e+17, 1.288744262932095e+17, 1.288744262972719e+17, 1.288744263013345e+17, 1.288744263052407e+17, 1.288744263093033e+17, 1.288744263132095e+17, 1.288744263172721e+17, 1.288744263213345e+17, 1.288744263252407e+17, 1.288744263293033e+17, 1.288744263332095e+17, 1.288744263372719e+17, 1.288744263413345e+17, 1.288744263452407e+17, 1.288744263493033e+17, 1.288744263532095e+17, 1.288744263572721e+17, 1.288744263613345e+17, 1.288744263652408e+17, 1.288744263693033e+17, 1.288744263732095e+17, 1.288744263772721e+17, 1.288744263813344e+17, 1.288744263852407e+17, 1.288744263893033e+17, 1.288744263932095e+17, 1.288744263972721e+17, 1.288744264013345e+17, 1.288744264052408e+17, 1.288744264093032e+17, 1.288744264132095e+17, 1.288744264172721e+17, 1.288744264213344e+17, 1.288744264252408e+17, 1.288744264293032e+17, 1.288744264332095e+17, 1.288744264372719e+17, 1.288744264413345e+17, 1.288744264452408e+17, 1.288744264493032e+17, 1.288744264532096e+17, 1.288744264572719e+17, 1.288744264613345e+17, 1.288744264652407e+17, 1.288744264693032e+17, 1.288744264732095e+17, 1.288744264772719e+17, 1.288744264813345e+17, 1.288744264852407e+17, 1.288744264893033e+17, 1.288744264932095e+17, 1.288744264972719e+17, 1.288744265013345e+17, 1.288744265052407e+17, 1.288744265093032e+17, 1.288744265132095e+17, 1.288744265172719e+17, 1.288744265213345e+17, 1.288744265252407e+17, 1.288744265293033e+17, 1.288744265332095e+17, 1.288744265372719e+17, 1.288744265413345e+17, 1.288744265452407e+17, 1.288744265493033e+17, 1.288744265532095e+17, 1.288744265572719e+17, 1.288744265613345e+17, 1.288744265652407e+17, 1.288744265693033e+17, 1.288744265732095e+17, 1.288744265772721e+17, 1.288744265813345e+17, 1.288744265852407e+17, 1.288744265893033e+17, 1.288744265932095e+17, 1.288744265972719e+17, 1.288744266013345e+17, 1.288744266052407e+17, 1.288744266093033e+17, 1.288744266132095e+17, 1.288744266172721e+17, 1.288744266213345e+17, 1.288744266252408e+17, 1.288744266293033e+17, 1.288744266332095e+17, 1.288744266372721e+17, 1.288744266413344e+17, 1.288744266452407e+17, 1.288744266493033e+17, 1.288744266532095e+17, 1.288744266572721e+17, 1.288744266613345e+17, 1.288744266652408e+17, 1.288744266693032e+17, 1.288744266732095e+17, 1.288744266772721e+17, 1.288744266813344e+17, 1.288744266852408e+17, 1.288744266893032e+17, 1.288744266932095e+17, 1.288744266972719e+17, 1.288744267013345e+17, 1.288744267052408e+17, 1.288744267093032e+17, 1.288744267132096e+17, 1.288744267172719e+17, 1.288744267213345e+17, 1.288744267252407e+17, 1.288744267293032e+17, 1.288744267332095e+17, 1.288744267372719e+17, 1.288744267413345e+17, 1.288744267452407e+17, 1.288744267493033e+17, 1.288744267532095e+17},
			             {1.288744306213345e+17, 1.288744306252407e+17, 1.288744306293033e+17, 1.288744306332095e+17, 1.288744306372719e+17, 1.288744306413345e+17, 1.288744306452407e+17, 1.288744306493033e+17, 1.288744306532095e+17, 1.288744306572721e+17, 1.288744306613345e+17, 1.288744306652407e+17, 1.288744306693033e+17, 1.288744306732095e+17, 1.288744306772721e+17, 1.288744306813345e+17, 1.288744306852407e+17, 1.288744306893033e+17, 1.288744306932095e+17, 1.288744306972721e+17, 1.288744307013345e+17, 1.288744307052408e+17, 1.288744307093033e+17, 1.288744307132095e+17, 1.288744307172721e+17, 1.288744307213344e+17, 1.288744307252407e+17, 1.288744307293033e+17, 1.288744307332095e+17, 1.288744307372721e+17, 1.288744307413345e+17, 1.288744307452408e+17, 1.288744307493032e+17, 1.288744307532095e+17, 1.288744307572721e+17, 1.288744307613344e+17, 1.288744307652408e+17, 1.288744307693032e+17, 1.288744307732095e+17, 1.288744307772719e+17, 1.288744307813345e+17, 1.288744307852408e+17, 1.288744307893032e+17, 1.288744307932096e+17, 1.288744307972719e+17, 1.288744308013345e+17, 1.288744308052407e+17, 1.288744308093032e+17, 1.288744308132095e+17, 1.288744308172719e+17, 1.288744308213345e+17, 1.288744308252407e+17, 1.288744308293033e+17, 1.288744308332095e+17, 1.288744308372719e+17, 1.288744308413345e+17},
			             {1.288744320652407e+17, 1.288744320693032e+17, 1.288744320732095e+17, 1.288744320772719e+17, 1.288744320813345e+17, 1.288744320852407e+17, 1.288744320893033e+17, 1.288744320932095e+17, 1.288744320972719e+17, 1.288744321013345e+17, 1.288744321052407e+17, 1.288744321093032e+17, 1.288744321132095e+17, 1.288744321172719e+17, 1.288744321213345e+17, 1.288744321252407e+17, 1.288744321293033e+17, 1.288744321332095e+17, 1.288744321372719e+17, 1.288744321413345e+17, 1.288744321452407e+17, 1.288744321493033e+17, 1.288744321532095e+17, 1.288744321572719e+17, 1.288744321613345e+17, 1.288744321652407e+17, 1.288744321693033e+17, 1.288744321732095e+17, 1.288744321772721e+17, 1.288744321813345e+17, 1.288744321852407e+17, 1.288744321893033e+17, 1.288744321932095e+17, 1.288744321972719e+17, 1.288744322013345e+17, 1.288744322052407e+17, 1.288744322093033e+17, 1.288744322132095e+17, 1.288744322172721e+17, 1.288744322213345e+17, 1.288744322252408e+17, 1.288744322293033e+17, 1.288744322332095e+17, 1.288744322372721e+17, 1.288744322413344e+17, 1.288744322452407e+17, 1.288744322493033e+17, 1.288744322532095e+17, 1.288744322572721e+17, 1.288744322613345e+17, 1.288744322652408e+17, 1.288744322693032e+17, 1.288744322732095e+17, 1.288744322772721e+17, 1.288744322813344e+17, 1.288744322852408e+17, 1.288744322893032e+17, 1.288744322932095e+17, 1.288744322972719e+17, 1.288744323013345e+17, 1.288744323052408e+17, 1.288744323093032e+17, 1.288744323132096e+17, 1.288744323172719e+17, 1.288744323213345e+17, 1.288744323252407e+17, 1.288744323293032e+17, 1.288744323332095e+17, 1.288744323372719e+17, 1.288744323413345e+17, 1.288744323452407e+17, 1.288744323493033e+17, 1.288744323532095e+17, 1.288744323572719e+17, 1.288744323613345e+17, 1.288744323652407e+17, 1.288744323693032e+17, 1.288744323732095e+17, 1.288744323772719e+17, 1.288744323813345e+17, 1.288744323852407e+17, 1.288744323893033e+17, 1.288744323932095e+17, 1.288744323972721e+17, 1.288744324013345e+17, 1.288744324052407e+17, 1.288744324093033e+17, 1.288744324132095e+17},
			             {1.288744231693032e+17, 1.288744231732095e+17, 1.288744231772719e+17, 1.288744231813345e+17, 1.288744231852407e+17, 1.288744231893033e+17, 1.288744231932095e+17},
			             {1.288744233813344e+17, 1.288744233852408e+17, 1.288744233893032e+17, 1.288744233932095e+17, 1.288744233972719e+17, 1.288744234013345e+17, 1.288744234052407e+17, 1.288744234093033e+17, 1.288744234132096e+17, 1.288744234172719e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
