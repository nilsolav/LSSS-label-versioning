netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 1;
			channels = 1;
			categories = 1;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0;
			max_depth =  246.3;
			start_time = 127825457244399488;
			end_time = 127825505795759488;
			region_id = 1;
			region_name = "Layer1";
			region_provenance = "LSSS";
			region_comment = "";
			region_category_names = "0";
			region_category_proportions = 1.0;
			region_category_ids = 1;
			region_type = analysis;
			channel_names = "";
			region_channels = 1;
			mask_times = {1.278254572443995e+17, 1.278254572543995e+17, 1.278254572643995e+17, 1.278254572743995e+17, 1.278254572843995e+17, 1.278254572943996e+17, 1.278254573043995e+17, 1.278254573143995e+17, 1.278254573243995e+17, 1.278254573343995e+17, 1.278254573443995e+17, 1.278254573543995e+17, 1.278254573643995e+17, 1.278254573743995e+17, 1.278254573843995e+17, 1.278254573943995e+17, 1.278254574043995e+17, 1.278254574143995e+17, 1.278254574243995e+17, 1.278254574343995e+17, 1.278254574443996e+17, 1.278254574543995e+17, 1.278254574643995e+17, 1.278254574743995e+17, 1.278254574843995e+17, 1.278254574943995e+17, 1.278254575043995e+17, 1.278254575143995e+17, 1.278254575243995e+17, 1.278254575343995e+17, 1.278254575443995e+17, 1.278254575543996e+17, 1.278254575643995e+17, 1.278254575743995e+17, 1.278254575843995e+17, 1.278254575943995e+17, 1.278254576043995e+17, 1.278254576143995e+17, 1.278254576243995e+17, 1.278254576343995e+17, 1.278254576443995e+17, 1.278254576543995e+17, 1.278254576643996e+17, 1.278254576743995e+17, 1.278254576843995e+17, 1.278254576943995e+17, 1.278254577043996e+17, 1.278254577143995e+17, 1.278254577243995e+17, 1.278254577343995e+17, 1.278254577443995e+17, 1.278254577543995e+17, 1.278254577643995e+17, 1.278254577743995e+17, 1.278254577843995e+17, 1.278254577943995e+17, 1.278254578043995e+17, 1.278254578143996e+17, 1.278254578243995e+17, 1.278254578343995e+17, 1.278254578443995e+17, 1.278254578543995e+17, 1.278254578643995e+17, 1.278254578743995e+17, 1.278254578843995e+17, 1.278254578943995e+17, 1.278254579043995e+17, 1.278254579143995e+17, 1.278254579243996e+17, 1.278254579343995e+17, 1.278254579443995e+17, 1.278254579543995e+17, 1.278254579643996e+17, 1.278254579743995e+17, 1.278254579843995e+17, 1.278254579943995e+17, 1.278254580043995e+17, 1.278254580143995e+17, 1.278254580243995e+17, 1.278254580343995e+17, 1.278254580443995e+17, 1.278254580543995e+17, 1.278254580643995e+17, 1.278254580743996e+17, 1.278254580843995e+17, 1.278254580943995e+17, 1.278254581043995e+17, 1.278254581143995e+17, 1.278254581243995e+17, 1.278254581343995e+17, 1.278254581443995e+17, 1.278254581543995e+17, 1.278254581643995e+17, 1.278254581743995e+17, 1.278254581843996e+17, 1.278254581943995e+17, 1.278254582043995e+17, 1.278254582143995e+17, 1.278254582243995e+17, 1.278254582343995e+17, 1.278254582443995e+17, 1.278254582543995e+17, 1.278254582643995e+17, 1.278254582743995e+17, 1.278254582843995e+17, 1.278254582943995e+17, 1.278254583043995e+17, 1.278254583143995e+17, 1.278254583243995e+17, 1.278254583343996e+17, 1.278254583443995e+17, 1.278254583543995e+17, 1.278254583643995e+17, 1.278254583743995e+17, 1.278254583843995e+17, 1.278254583943995e+17, 1.278254584043995e+17, 1.278254584143995e+17, 1.278254584243995e+17, 1.278254584343995e+17, 1.278254584443996e+17, 1.278254584543995e+17, 1.278254584643995e+17, 1.278254584743995e+17, 1.278254584843995e+17, 1.278254584943995e+17, 1.278254585043995e+17, 1.278254585143995e+17, 1.278254585243995e+17, 1.278254585343995e+17, 1.278254585443995e+17, 1.278254585543995e+17, 1.278254585643995e+17, 1.278254585743995e+17, 1.278254585843995e+17, 1.278254585943996e+17, 1.278254586043995e+17, 1.278254586143995e+17, 1.278254586243995e+17, 1.278254586343995e+17, 1.278254586443995e+17, 1.278254586543995e+17, 1.278254586643995e+17, 1.278254586743995e+17, 1.278254586843995e+17, 1.278254586943995e+17, 1.278254587043996e+17, 1.278254587143995e+17, 1.278254587243995e+17, 1.278254587343995e+17, 1.278254587443995e+17, 1.278254587543995e+17, 1.278254587643995e+17, 1.278254587743995e+17, 1.278254587843995e+17, 1.278254587943995e+17, 1.278254588043995e+17, 1.278254588143996e+17, 1.278254588243995e+17, 1.278254588343995e+17, 1.278254588443995e+17, 1.278254588543996e+17, 1.278254588643995e+17, 1.278254588743995e+17, 1.278254588843995e+17, 1.278254588943995e+17, 1.278254589043995e+17, 1.278254589143995e+17, 1.278254589243995e+17, 1.278254589343995e+17, 1.278254589443995e+17, 1.278254589543995e+17, 1.278254589643996e+17, 1.278254589743995e+17, 1.278254589843995e+17, 1.278254589943995e+17, 1.278254590043995e+17, 1.278254590143995e+17, 1.278254590243995e+17, 1.278254590343995e+17, 1.278254590443995e+17, 1.278254590543995e+17, 1.278254590643995e+17, 1.278254590743996e+17, 1.278254590843995e+17, 1.278254590943995e+17, 1.278254591043995e+17, 1.278254591143996e+17, 1.278254591243995e+17, 1.278254591343995e+17, 1.278254591443995e+17, 1.278254591543995e+17, 1.278254591643995e+17, 1.278254591743995e+17, 1.278254591843995e+17, 1.278254591943995e+17, 1.278254592043995e+17, 1.278254592143995e+17, 1.278254592243996e+17, 1.278254592343995e+17, 1.278254592443995e+17, 1.278254592543995e+17, 1.278254592643995e+17, 1.278254592743995e+17, 1.278254592843995e+17, 1.278254592943995e+17, 1.278254593043995e+17, 1.278254593143995e+17, 1.278254593243995e+17, 1.278254593343996e+17, 1.278254593443995e+17, 1.278254593543995e+17, 1.278254593643995e+17, 1.278254593743995e+17, 1.278254593843995e+17, 1.278254593943995e+17, 1.278254594043995e+17, 1.278254594143995e+17, 1.278254594243995e+17, 1.278254594343995e+17, 1.278254594443995e+17, 1.278254594543995e+17, 1.278254594643995e+17, 1.278254594743995e+17, 1.278254594843996e+17, 1.278254594943995e+17, 1.278254595043995e+17, 1.278254595143995e+17, 1.278254595243995e+17, 1.278254595343995e+17, 1.278254595443995e+17, 1.278254595543995e+17, 1.278254595643995e+17, 1.278254595743995e+17, 1.278254595843995e+17, 1.278254595943996e+17, 1.278254596043995e+17, 1.278254596143995e+17, 1.278254596243995e+17, 1.278254596343995e+17, 1.278254596443995e+17, 1.278254596543995e+17, 1.278254596643995e+17, 1.278254596743995e+17, 1.278254596843995e+17, 1.278254596943995e+17, 1.278254597043996e+17, 1.278254597143995e+17, 1.278254597243995e+17, 1.278254597343995e+17, 1.278254597443996e+17, 1.278254597543995e+17, 1.278254597643995e+17, 1.278254597743995e+17, 1.278254597843995e+17, 1.278254597943995e+17, 1.278254598043995e+17, 1.278254598143995e+17, 1.278254598243995e+17, 1.278254598343995e+17, 1.278254598443995e+17, 1.278254598543996e+17, 1.278254598643995e+17, 1.278254598743995e+17, 1.278254598843995e+17, 1.278254598943995e+17, 1.278254599043995e+17, 1.278254599143995e+17, 1.278254599243995e+17, 1.278254599343995e+17, 1.278254599443995e+17, 1.278254599543995e+17, 1.278254599643996e+17, 1.278254599743995e+17, 1.278254599843995e+17, 1.278254599943995e+17, 1.278254600043996e+17, 1.278254600143995e+17, 1.278254600243995e+17, 1.278254600343995e+17, 1.278254600443995e+17, 1.278254600543995e+17, 1.278254600643995e+17, 1.278254600743995e+17, 1.278254600843995e+17, 1.278254600943995e+17, 1.278254601043995e+17, 1.278254601143996e+17, 1.278254601243995e+17, 1.278254601343995e+17, 1.278254601443995e+17, 1.278254601543995e+17, 1.278254601643995e+17, 1.278254601743995e+17, 1.278254601843995e+17, 1.278254601943995e+17, 1.278254602043995e+17, 1.278254602143995e+17, 1.278254602243996e+17, 1.278254602343995e+17, 1.278254602443995e+17, 1.278254602543995e+17, 1.278254602643995e+17, 1.278254602743995e+17, 1.278254602843995e+17, 1.278254602943995e+17, 1.278254603043995e+17, 1.278254603143995e+17, 1.278254603243995e+17, 1.278254603343995e+17, 1.278254603443995e+17, 1.278254603543995e+17, 1.278254603643995e+17, 1.278254603743996e+17, 1.278254603843995e+17, 1.278254603943995e+17, 1.278254604043995e+17, 1.278254604143995e+17, 1.278254604243995e+17, 1.278254604343995e+17, 1.278254604443995e+17, 1.278254604543995e+17, 1.278254604643995e+17, 1.278254604743995e+17, 1.278254604843996e+17, 1.278254604943995e+17, 1.278254605043995e+17, 1.278254605143995e+17, 1.278254605243995e+17, 1.278254605343995e+17, 1.278254605443995e+17, 1.278254605543995e+17, 1.278254605643995e+17, 1.278254605743995e+17, 1.278254605843995e+17, 1.278254605943996e+17, 1.278254606043995e+17, 1.278254606143995e+17, 1.278254606243995e+17, 1.278254606343996e+17, 1.278254606443995e+17, 1.278254606543995e+17, 1.278254606643995e+17, 1.278254606743995e+17, 1.278254606843995e+17, 1.278254606943995e+17, 1.278254607043995e+17, 1.278254607143995e+17, 1.278254607243995e+17, 1.278254607343995e+17, 1.278254607443996e+17, 1.278254607543995e+17, 1.278254607643995e+17, 1.278254607743995e+17, 1.278254607843995e+17, 1.278254607943995e+17, 1.278254608043995e+17, 1.278254608143995e+17, 1.278254608243995e+17, 1.278254608343995e+17, 1.278254608443995e+17, 1.278254608543996e+17, 1.278254608643995e+17, 1.278254608743995e+17, 1.278254608843995e+17, 1.278254608943996e+17, 1.278254609043995e+17, 1.278254609143995e+17, 1.278254609243995e+17, 1.278254609343995e+17, 1.278254609443995e+17, 1.278254609543995e+17, 1.278254609643995e+17, 1.278254609743995e+17, 1.278254609843995e+17, 1.278254609943995e+17, 1.278254610043996e+17, 1.278254610143995e+17, 1.278254610243995e+17, 1.278254610343995e+17, 1.278254610443995e+17, 1.278254610543995e+17, 1.278254610643995e+17, 1.278254610743995e+17, 1.278254610843995e+17, 1.278254610943995e+17, 1.278254611043995e+17, 1.278254611143996e+17, 1.278254611243995e+17, 1.278254611343995e+17, 1.278254611443995e+17, 1.278254611543995e+17, 1.278254611643995e+17, 1.278254611743995e+17, 1.278254611843995e+17, 1.278254611943995e+17, 1.278254612043995e+17, 1.278254612143995e+17, 1.278254612243995e+17, 1.278254612343995e+17, 1.278254612443995e+17, 1.278254612543995e+17, 1.278254612643996e+17, 1.278254612743995e+17, 1.278254612843995e+17, 1.278254612943995e+17, 1.278254613043995e+17, 1.278254613143995e+17, 1.278254613243995e+17, 1.278254613343995e+17, 1.278254613443995e+17, 1.278254613543995e+17, 1.278254613643995e+17, 1.278254613743996e+17, 1.278254613843995e+17, 1.278254613943995e+17, 1.278254614043995e+17, 1.278254614143995e+17, 1.278254614243995e+17, 1.278254614343995e+17, 1.278254614443995e+17, 1.278254614543995e+17, 1.278254614643995e+17, 1.278254614743995e+17, 1.278254614843996e+17, 1.278254614943995e+17, 1.278254615043995e+17, 1.278254615143995e+17, 1.278254615243996e+17, 1.278254615343995e+17, 1.278254615443995e+17, 1.278254615543995e+17, 1.278254615643995e+17, 1.278254615743995e+17, 1.278254615843995e+17, 1.278254615943995e+17, 1.278254616043995e+17, 1.278254616143995e+17, 1.278254616243995e+17, 1.278254616343996e+17, 1.278254616443995e+17, 1.278254616543995e+17, 1.278254616643995e+17, 1.278254616743995e+17, 1.278254616843995e+17, 1.278254616943995e+17, 1.278254617043995e+17, 1.278254617143995e+17, 1.278254617243995e+17, 1.278254617343995e+17, 1.278254617443996e+17, 1.278254617543995e+17, 1.278254617643995e+17, 1.278254617743995e+17, 1.278254617843996e+17, 1.278254617943995e+17, 1.278254618043995e+17, 1.278254618143995e+17, 1.278254618243995e+17, 1.278254618343995e+17, 1.278254618443995e+17, 1.278254618543995e+17, 1.278254618643995e+17, 1.278254618743995e+17, 1.278254618843995e+17, 1.278254618943996e+17, 1.278254619043995e+17, 1.278254619143995e+17, 1.278254619243995e+17, 1.278254619343995e+17, 1.278254619443995e+17, 1.278254619543995e+17, 1.278254619643995e+17, 1.278254619743995e+17, 1.278254619843995e+17, 1.278254619943995e+17, 1.278254620043996e+17, 1.278254620143995e+17, 1.278254620243995e+17, 1.278254620343995e+17, 1.278254620443996e+17, 1.278254620543995e+17, 1.278254620643995e+17, 1.278254620743995e+17, 1.278254620843995e+17, 1.278254620943995e+17, 1.278254621043995e+17, 1.278254621143995e+17, 1.278254621243995e+17, 1.278254621343995e+17, 1.278254621443995e+17, 1.278254621543996e+17, 1.278254621643995e+17, 1.278254621743995e+17, 1.278254621843995e+17, 1.278254621943995e+17, 1.278254622043995e+17, 1.278254622143995e+17, 1.278254622243995e+17, 1.278254622343995e+17, 1.278254622443995e+17, 1.278254622543995e+17, 1.278254622643996e+17, 1.278254622743995e+17, 1.278254622843995e+17, 1.278254622943995e+17, 1.278254623043995e+17, 1.278254623143995e+17, 1.278254623243995e+17, 1.278254623343995e+17, 1.278254623443995e+17, 1.278254623543995e+17, 1.278254623643995e+17, 1.278254623743995e+17, 1.278254623843995e+17, 1.278254623943995e+17, 1.278254624043995e+17, 1.278254624143996e+17, 1.278254624243995e+17, 1.278254624343995e+17, 1.278254624443995e+17, 1.278254624543995e+17, 1.278254624643995e+17, 1.278254624743995e+17, 1.278254624843995e+17, 1.278254624943995e+17, 1.278254625043995e+17, 1.278254625143995e+17, 1.278254625243996e+17, 1.278254625343995e+17, 1.278254625443995e+17, 1.278254625543995e+17, 1.278254625643995e+17, 1.278254625743995e+17, 1.278254625843995e+17, 1.278254625943995e+17, 1.278254626043995e+17, 1.278254626143995e+17, 1.278254626243995e+17, 1.278254626343996e+17, 1.278254626443995e+17, 1.278254626543995e+17, 1.278254626643995e+17, 1.278254626743996e+17, 1.278254626843995e+17, 1.278254626943995e+17, 1.278254627043995e+17, 1.278254627143995e+17, 1.278254627243995e+17, 1.278254627343995e+17, 1.278254627443995e+17, 1.278254627543995e+17, 1.278254627643995e+17, 1.278254627743995e+17, 1.278254627843996e+17, 1.278254627943995e+17, 1.278254628043995e+17, 1.278254628143995e+17, 1.278254628243995e+17, 1.278254628343995e+17, 1.278254628443995e+17, 1.278254628543995e+17, 1.278254628643995e+17, 1.278254628743995e+17, 1.278254628843995e+17, 1.278254628943996e+17, 1.278254629043995e+17, 1.278254629143995e+17, 1.278254629243995e+17, 1.278254629343996e+17, 1.278254629443995e+17, 1.278254629543995e+17, 1.278254629643995e+17, 1.278254629743995e+17, 1.278254629843995e+17, 1.278254629943995e+17, 1.278254630043995e+17, 1.278254630143995e+17, 1.278254630243995e+17, 1.278254630343995e+17, 1.278254630443996e+17, 1.278254630543995e+17, 1.278254630643995e+17, 1.278254630743995e+17, 1.278254630843995e+17, 1.278254630943995e+17, 1.278254631043995e+17, 1.278254631143995e+17, 1.278254631243995e+17, 1.278254631343995e+17, 1.278254631443995e+17, 1.278254631543996e+17, 1.278254631643995e+17, 1.278254631743995e+17, 1.278254631843995e+17, 1.278254631943995e+17, 1.278254632043995e+17, 1.278254632143995e+17, 1.278254632243995e+17, 1.278254632343995e+17, 1.278254632443995e+17, 1.278254632543995e+17, 1.278254632643995e+17, 1.278254632743995e+17, 1.278254632843995e+17, 1.278254632943995e+17, 1.278254633043996e+17, 1.278254633143995e+17, 1.278254633243995e+17, 1.278254633343995e+17, 1.278254633443995e+17, 1.278254633543995e+17, 1.278254633643995e+17, 1.278254633743995e+17, 1.278254633843995e+17, 1.278254633943995e+17, 1.278254634043995e+17, 1.278254634143996e+17, 1.278254634243995e+17, 1.278254634343995e+17, 1.278254634443995e+17, 1.278254634543995e+17, 1.278254634643995e+17, 1.278254634743995e+17, 1.278254634843995e+17, 1.278254634943995e+17, 1.278254635043995e+17, 1.278254635143995e+17, 1.278254635243996e+17, 1.278254635343995e+17, 1.278254635443995e+17, 1.278254635543995e+17, 1.278254635643996e+17, 1.278254635743995e+17, 1.278254635843995e+17, 1.278254635943995e+17, 1.278254636043995e+17, 1.278254636143995e+17, 1.278254636243995e+17, 1.278254636343995e+17, 1.278254636443995e+17, 1.278254636543995e+17, 1.278254636643995e+17, 1.278254636743996e+17, 1.278254636843995e+17, 1.278254636943995e+17, 1.278254637043995e+17, 1.278254637143995e+17, 1.278254637243995e+17, 1.278254637343995e+17, 1.278254637443995e+17, 1.278254637543995e+17, 1.278254637643995e+17, 1.278254637743995e+17, 1.278254637843996e+17, 1.278254637943995e+17, 1.278254638043995e+17, 1.278254638143995e+17, 1.278254638243996e+17, 1.278254638343995e+17, 1.278254638443995e+17, 1.278254638543995e+17, 1.278254638643995e+17, 1.278254638743995e+17, 1.278254638843995e+17, 1.278254638943995e+17, 1.278254639043995e+17, 1.278254639143995e+17, 1.278254639243995e+17, 1.278254639343996e+17, 1.278254639443995e+17, 1.278254639543995e+17, 1.278254639643995e+17, 1.278254639743995e+17, 1.278254639843995e+17, 1.278254639943995e+17, 1.278254640043995e+17, 1.278254640143995e+17, 1.278254640243995e+17, 1.278254640343995e+17, 1.278254640443996e+17, 1.278254640543995e+17, 1.278254640643995e+17, 1.278254640743995e+17, 1.278254640843995e+17, 1.278254640943995e+17, 1.278254641043995e+17, 1.278254641143995e+17, 1.278254641243995e+17, 1.278254641343995e+17, 1.278254641443995e+17, 1.278254641543995e+17, 1.278254641643995e+17, 1.278254641743995e+17, 1.278254641843995e+17, 1.278254641943996e+17, 1.278254642043995e+17, 1.278254642143995e+17, 1.278254642243995e+17, 1.278254642343995e+17, 1.278254642443995e+17, 1.278254642543995e+17, 1.278254642643995e+17, 1.278254642743995e+17, 1.278254642843995e+17, 1.278254642943995e+17, 1.278254643043996e+17, 1.278254643143995e+17, 1.278254643243995e+17, 1.278254643343995e+17, 1.278254643443995e+17, 1.278254643543995e+17, 1.278254643643995e+17, 1.278254643743995e+17, 1.278254643843995e+17, 1.278254643943995e+17, 1.278254644043995e+17, 1.278254644143996e+17, 1.278254644243995e+17, 1.278254644343995e+17, 1.278254644443995e+17, 1.278254644543996e+17, 1.278254644643995e+17, 1.278254644743995e+17, 1.278254644843995e+17, 1.278254644943995e+17, 1.278254645043995e+17, 1.278254645143995e+17, 1.278254645243995e+17, 1.278254645343995e+17, 1.278254645443995e+17, 1.278254645543995e+17, 1.278254645643996e+17, 1.278254645743995e+17, 1.278254645843995e+17, 1.278254645943995e+17, 1.278254646043995e+17, 1.278254646143995e+17, 1.278254646243995e+17, 1.278254646343995e+17, 1.278254646443995e+17, 1.278254646543995e+17, 1.278254646643995e+17, 1.278254646743996e+17, 1.278254646843995e+17, 1.278254646943995e+17, 1.278254647043995e+17, 1.278254647143996e+17, 1.278254647243995e+17, 1.278254647343995e+17, 1.278254647443995e+17, 1.278254647543995e+17, 1.278254647643995e+17, 1.278254647743995e+17, 1.278254647843995e+17, 1.278254647943995e+17, 1.278254648043995e+17, 1.278254648143995e+17, 1.278254648243996e+17, 1.278254648343995e+17, 1.278254648443995e+17, 1.278254648543995e+17, 1.278254648643995e+17, 1.278254648743995e+17, 1.278254648843995e+17, 1.278254648943995e+17, 1.278254649043995e+17, 1.278254649143995e+17, 1.278254649243995e+17, 1.278254649343996e+17, 1.278254649443995e+17, 1.278254649543995e+17, 1.278254649643995e+17, 1.278254649743995e+17, 1.278254649843995e+17, 1.278254649943995e+17, 1.278254650043995e+17, 1.278254650143995e+17, 1.278254650243995e+17, 1.278254650343995e+17, 1.278254650443995e+17, 1.278254650543995e+17, 1.278254650643995e+17, 1.278254650743995e+17, 1.278254650843996e+17, 1.278254650943995e+17, 1.278254651043995e+17, 1.278254651143995e+17, 1.278254651243995e+17, 1.278254651343995e+17, 1.278254651443995e+17, 1.278254651543995e+17, 1.278254651643995e+17, 1.278254651743995e+17, 1.278254651843995e+17, 1.278254651943996e+17, 1.278254652043995e+17, 1.278254652143995e+17, 1.278254652243995e+17, 1.278254652343995e+17, 1.278254652443995e+17, 1.278254652543995e+17, 1.278254652643995e+17, 1.278254652743995e+17, 1.278254652843995e+17, 1.278254652943995e+17, 1.278254653043995e+17, 1.278254653143995e+17, 1.278254653243995e+17, 1.278254653343995e+17, 1.278254653443996e+17, 1.278254653543995e+17, 1.278254653643995e+17, 1.278254653743995e+17, 1.278254653843995e+17, 1.278254653943995e+17, 1.278254654043995e+17, 1.278254654143995e+17, 1.278254654243995e+17, 1.278254654343995e+17, 1.278254654443995e+17, 1.278254654543996e+17, 1.278254654643995e+17, 1.278254654743995e+17, 1.278254654843995e+17, 1.278254654943995e+17, 1.278254655043995e+17, 1.278254655143995e+17, 1.278254655243995e+17, 1.278254655343995e+17, 1.278254655443995e+17, 1.278254655543995e+17, 1.278254655643996e+17, 1.278254655743995e+17, 1.278254655843995e+17, 1.278254655943995e+17, 1.278254656043996e+17, 1.278254656143995e+17, 1.278254656243995e+17, 1.278254656343995e+17, 1.278254656443995e+17, 1.278254656543995e+17, 1.278254656643995e+17, 1.278254656743995e+17, 1.278254656843995e+17, 1.278254656943995e+17, 1.278254657043995e+17, 1.278254657143996e+17, 1.278254657243995e+17, 1.278254657343995e+17, 1.278254657443995e+17, 1.278254657543995e+17, 1.278254657643995e+17, 1.278254657743995e+17, 1.278254657843995e+17, 1.278254657943995e+17, 1.278254658043995e+17, 1.278254658143995e+17, 1.278254658243996e+17, 1.278254658343995e+17, 1.278254658443995e+17, 1.278254658543995e+17, 1.278254658643996e+17, 1.278254658743995e+17, 1.278254658843995e+17, 1.278254658943995e+17, 1.278254659043995e+17, 1.278254659143995e+17, 1.278254659243995e+17, 1.278254659343995e+17, 1.278254659443995e+17, 1.278254659543995e+17, 1.278254659643995e+17, 1.278254659743996e+17, 1.278254659843995e+17, 1.278254659943995e+17, 1.278254660043995e+17, 1.278254660143995e+17, 1.278254660243995e+17, 1.278254660343995e+17, 1.278254660443995e+17, 1.278254660543995e+17, 1.278254660643995e+17, 1.278254660743995e+17, 1.278254660843996e+17, 1.278254660943995e+17, 1.278254661043995e+17, 1.278254661143995e+17, 1.278254661243995e+17, 1.278254661343995e+17, 1.278254661443995e+17, 1.278254661543995e+17, 1.278254661643995e+17, 1.278254661743995e+17, 1.278254661843995e+17, 1.278254661943995e+17, 1.278254662043995e+17, 1.278254662143995e+17, 1.278254662243995e+17, 1.278254662343996e+17, 1.278254662443995e+17, 1.278254662543995e+17, 1.278254662643995e+17, 1.278254662743995e+17, 1.278254662843995e+17, 1.278254662943995e+17, 1.278254663043995e+17, 1.278254663143995e+17, 1.278254663243995e+17, 1.278254663343995e+17, 1.278254663443996e+17, 1.278254663543995e+17, 1.278254663643995e+17, 1.278254663743995e+17, 1.278254663843995e+17, 1.278254663943995e+17, 1.278254664043995e+17, 1.278254664143995e+17, 1.278254664243995e+17, 1.278254664343995e+17, 1.278254664443995e+17, 1.278254664543996e+17, 1.278254664643995e+17, 1.278254664743995e+17, 1.278254664843995e+17, 1.278254664943996e+17, 1.278254665043995e+17, 1.278254665143995e+17, 1.278254665243995e+17, 1.278254665343995e+17, 1.278254665443995e+17, 1.278254665543995e+17, 1.278254665643995e+17, 1.278254665743995e+17, 1.278254665843995e+17, 1.278254665943995e+17, 1.278254666043996e+17, 1.278254666143995e+17, 1.278254666243995e+17, 1.278254666343995e+17, 1.278254666443995e+17, 1.278254666543995e+17, 1.278254666643995e+17, 1.278254666743995e+17, 1.278254666843995e+17, 1.278254666943995e+17, 1.278254667043995e+17, 1.278254667143996e+17, 1.278254667243995e+17, 1.278254667343995e+17, 1.278254667443995e+17, 1.278254667543996e+17, 1.278254667643995e+17, 1.278254667743995e+17, 1.278254667843995e+17, 1.278254667943995e+17, 1.278254668043995e+17, 1.278254668143995e+17, 1.278254668243995e+17, 1.278254668343995e+17, 1.278254668443995e+17, 1.278254668543995e+17, 1.278254668643996e+17, 1.278254668743995e+17, 1.278254668843995e+17, 1.278254668943995e+17, 1.278254669043995e+17, 1.278254669143995e+17, 1.278254669243995e+17, 1.278254669343995e+17, 1.278254669443995e+17, 1.278254669543995e+17, 1.278254669643995e+17, 1.278254669743996e+17, 1.278254669843995e+17, 1.278254669943995e+17, 1.278254670043995e+17, 1.278254670143995e+17, 1.278254670243995e+17, 1.278254670343995e+17, 1.278254670443995e+17, 1.278254670543995e+17, 1.278254670643995e+17, 1.278254670743995e+17, 1.278254670843995e+17, 1.278254670943995e+17, 1.278254671043995e+17, 1.278254671143995e+17, 1.278254671243996e+17, 1.278254671343995e+17, 1.278254671443995e+17, 1.278254671543995e+17, 1.278254671643995e+17, 1.278254671743995e+17, 1.278254671843995e+17, 1.278254671943995e+17, 1.278254672043995e+17, 1.278254672143995e+17, 1.278254672243995e+17, 1.278254672343996e+17, 1.278254672443995e+17, 1.278254672543995e+17, 1.278254672643995e+17, 1.278254672743995e+17, 1.278254672843995e+17, 1.278254672943995e+17, 1.278254673043995e+17, 1.278254673143995e+17, 1.278254673243995e+17, 1.278254673343995e+17, 1.278254673443996e+17, 1.278254673543995e+17, 1.278254673643995e+17, 1.278254673743995e+17, 1.278254673843996e+17, 1.278254673943995e+17, 1.278254674043995e+17, 1.278254674143995e+17, 1.278254674243995e+17, 1.278254674343995e+17, 1.278254674443995e+17, 1.278254674543995e+17, 1.278254674643995e+17, 1.278254674743995e+17, 1.278254674843995e+17, 1.278254674943996e+17, 1.278254675043995e+17, 1.278254675143995e+17, 1.278254675243995e+17, 1.278254675343995e+17, 1.278254675443995e+17, 1.278254675543995e+17, 1.278254675643995e+17, 1.278254675743995e+17, 1.278254675843995e+17, 1.278254675943995e+17, 1.278254676043996e+17, 1.278254676143995e+17, 1.278254676243995e+17, 1.278254676343995e+17, 1.278254676443996e+17, 1.278254676543995e+17, 1.278254676643995e+17, 1.278254676743995e+17, 1.278254676843995e+17, 1.278254676943995e+17, 1.278254677043995e+17, 1.278254677143995e+17, 1.278254677243995e+17, 1.278254677343995e+17, 1.278254677443995e+17, 1.278254677543996e+17, 1.278254677643995e+17, 1.278254677743995e+17, 1.278254677843995e+17, 1.278254677943995e+17, 1.278254678043995e+17, 1.278254678143995e+17, 1.278254678243995e+17, 1.278254678343995e+17, 1.278254678443995e+17, 1.278254678543995e+17, 1.278254678643996e+17, 1.278254678743995e+17, 1.278254678843995e+17, 1.278254678943995e+17, 1.278254679043995e+17, 1.278254679143995e+17, 1.278254679243995e+17, 1.278254679343995e+17, 1.278254679443995e+17, 1.278254679543995e+17, 1.278254679643995e+17, 1.278254679743995e+17, 1.278254679843995e+17, 1.278254679943995e+17, 1.278254680043995e+17, 1.278254680143996e+17, 1.278254680243995e+17, 1.278254680343995e+17, 1.278254680443995e+17, 1.278254680543995e+17, 1.278254680643995e+17, 1.278254680743995e+17, 1.278254680843995e+17, 1.278254680943995e+17, 1.278254681043995e+17, 1.278254681143995e+17, 1.278254681243996e+17, 1.278254681343995e+17, 1.278254681443995e+17, 1.278254681543995e+17, 1.278254681643995e+17, 1.278254681743995e+17, 1.278254681843995e+17, 1.278254681943995e+17, 1.278254682043995e+17, 1.278254682143995e+17, 1.278254682243995e+17, 1.278254682343996e+17, 1.278254682443995e+17, 1.278254682543995e+17, 1.278254682643995e+17, 1.278254682743996e+17, 1.278254682843995e+17, 1.278254682943995e+17, 1.278254683043995e+17, 1.278254683143995e+17, 1.278254683243995e+17, 1.278254683343995e+17, 1.278254683443995e+17, 1.278254683543995e+17, 1.278254683643995e+17, 1.278254683743995e+17, 1.278254683843996e+17, 1.278254683943995e+17, 1.278254684043995e+17, 1.278254684143995e+17, 1.278254684243995e+17, 1.278254684343995e+17, 1.278254684443995e+17, 1.278254684543995e+17, 1.278254684643995e+17, 1.278254684743995e+17, 1.278254684843995e+17, 1.278254684943996e+17, 1.278254685043995e+17, 1.278254685143995e+17, 1.278254685243995e+17, 1.278254685343996e+17, 1.278254685443995e+17, 1.278254685543995e+17, 1.278254685643995e+17, 1.278254685743995e+17, 1.278254685843995e+17, 1.278254685943995e+17, 1.278254686043995e+17, 1.278254686143995e+17, 1.278254686243995e+17, 1.278254686343995e+17, 1.278254686443996e+17, 1.278254686543995e+17, 1.278254686643995e+17, 1.278254686743995e+17, 1.278254686843995e+17, 1.278254686943995e+17, 1.278254687043995e+17, 1.278254687143995e+17, 1.278254687243995e+17, 1.278254687343995e+17, 1.278254687443995e+17, 1.278254687543996e+17, 1.278254687643995e+17, 1.278254687743995e+17, 1.278254687843995e+17, 1.278254687943996e+17, 1.278254688043995e+17, 1.278254688143995e+17, 1.278254688243995e+17, 1.278254688343995e+17, 1.278254688443995e+17, 1.278254688543995e+17, 1.278254688643995e+17, 1.278254688743995e+17, 1.278254688843995e+17, 1.278254688943995e+17, 1.278254689043996e+17, 1.278254689143995e+17, 1.278254689243995e+17, 1.278254689343995e+17, 1.278254689443995e+17, 1.278254689543995e+17, 1.278254689643995e+17, 1.278254689743995e+17, 1.278254689843995e+17, 1.278254689943995e+17, 1.278254690043995e+17, 1.278254690143996e+17, 1.278254690243995e+17, 1.278254690343995e+17, 1.278254690443995e+17, 1.278254690543995e+17, 1.278254690643995e+17, 1.278254690743995e+17, 1.278254690843995e+17, 1.278254690943995e+17, 1.278254691043995e+17, 1.278254691143995e+17, 1.278254691243995e+17, 1.278254691343995e+17, 1.278254691443995e+17, 1.278254691543995e+17, 1.278254691643996e+17, 1.278254691743995e+17, 1.278254691843995e+17, 1.278254691943995e+17, 1.278254692043995e+17, 1.278254692143995e+17, 1.278254692243995e+17, 1.278254692343995e+17, 1.278254692443995e+17, 1.278254692543995e+17, 1.278254692643995e+17, 1.278254692743996e+17, 1.278254692843995e+17, 1.278254692943995e+17, 1.278254693043995e+17, 1.278254693143995e+17, 1.278254693243995e+17, 1.278254693343995e+17, 1.278254693443995e+17, 1.278254693543995e+17, 1.278254693643995e+17, 1.278254693743995e+17, 1.278254693843996e+17, 1.278254693943995e+17, 1.278254694043995e+17, 1.278254694143995e+17, 1.278254694243996e+17, 1.278254694343995e+17, 1.278254694443995e+17, 1.278254694543995e+17, 1.278254694643995e+17, 1.278254694743995e+17, 1.278254694843995e+17, 1.278254694943995e+17, 1.278254695043995e+17, 1.278254695143995e+17, 1.278254695243995e+17, 1.278254695343996e+17, 1.278254695443995e+17, 1.278254695543995e+17, 1.278254695643995e+17, 1.278254695743995e+17, 1.278254695843995e+17, 1.278254695943995e+17, 1.278254696043995e+17, 1.278254696143995e+17, 1.278254696243995e+17, 1.278254696343995e+17, 1.278254696443996e+17, 1.278254696543995e+17, 1.278254696643995e+17, 1.278254696743995e+17, 1.278254696843996e+17, 1.278254696943995e+17, 1.278254697043995e+17, 1.278254697143995e+17, 1.278254697243995e+17, 1.278254697343995e+17, 1.278254697443995e+17, 1.278254697543995e+17, 1.278254697643995e+17, 1.278254697743995e+17, 1.278254697843995e+17, 1.278254697943996e+17, 1.278254698043995e+17, 1.278254698143995e+17, 1.278254698243995e+17, 1.278254698343995e+17, 1.278254698443995e+17, 1.278254698543995e+17, 1.278254698643995e+17, 1.278254698743995e+17, 1.278254698843995e+17, 1.278254698943995e+17, 1.278254699043996e+17, 1.278254699143995e+17, 1.278254699243995e+17, 1.278254699343995e+17, 1.278254699443995e+17, 1.278254699543995e+17, 1.278254699643995e+17, 1.278254699743995e+17, 1.278254699843995e+17, 1.278254699943995e+17, 1.278254700043995e+17, 1.278254700143995e+17, 1.278254700243995e+17, 1.278254700343995e+17, 1.278254700443995e+17, 1.278254700543996e+17, 1.278254700643995e+17, 1.278254700743995e+17, 1.278254700843995e+17, 1.278254700943995e+17, 1.278254701043995e+17, 1.278254701143995e+17, 1.278254701243995e+17, 1.278254701343995e+17, 1.278254701443995e+17, 1.278254701543995e+17, 1.278254701643996e+17, 1.278254701743995e+17, 1.278254701843995e+17, 1.278254701943995e+17, 1.278254702043995e+17, 1.278254702143995e+17, 1.278254702243995e+17, 1.278254702343995e+17, 1.278254702443995e+17, 1.278254702543995e+17, 1.278254702643995e+17, 1.278254702743996e+17, 1.278254702843995e+17, 1.278254702943995e+17, 1.278254703043995e+17, 1.278254703143996e+17, 1.278254703243995e+17, 1.278254703343995e+17, 1.278254703443995e+17, 1.278254703543995e+17, 1.278254703643995e+17, 1.278254703743995e+17, 1.278254703843995e+17, 1.278254703943995e+17, 1.278254704043995e+17, 1.278254704143995e+17, 1.278254704243996e+17, 1.278254704343995e+17, 1.278254704443995e+17, 1.278254704543995e+17, 1.278254704643995e+17, 1.278254704743995e+17, 1.278254704843995e+17, 1.278254704943995e+17, 1.278254705043995e+17, 1.278254705143995e+17, 1.278254705243995e+17, 1.278254705343996e+17, 1.278254705443995e+17, 1.278254705543995e+17, 1.278254705643995e+17, 1.278254705743996e+17, 1.278254705843995e+17, 1.278254705943995e+17, 1.278254706043995e+17, 1.278254706143995e+17, 1.278254706243995e+17, 1.278254706343995e+17, 1.278254706443995e+17, 1.278254706543995e+17, 1.278254706643995e+17, 1.278254706743995e+17, 1.278254706843996e+17, 1.278254706943995e+17, 1.278254707043995e+17, 1.278254707143995e+17, 1.278254707243995e+17, 1.278254707343995e+17, 1.278254707443995e+17, 1.278254707543995e+17, 1.278254707643995e+17, 1.278254707743995e+17, 1.278254707843995e+17, 1.278254707943996e+17, 1.278254708043995e+17, 1.278254708143995e+17, 1.278254708243995e+17, 1.278254708343995e+17, 1.278254708443995e+17, 1.278254708543995e+17, 1.278254708643995e+17, 1.278254708743995e+17, 1.278254708843995e+17, 1.278254708943995e+17, 1.278254709043995e+17, 1.278254709143995e+17, 1.278254709243995e+17, 1.278254709343995e+17, 1.278254709443996e+17, 1.278254709543995e+17, 1.278254709643995e+17, 1.278254709743995e+17, 1.278254709843995e+17, 1.278254709943995e+17, 1.278254710043995e+17, 1.278254710143995e+17, 1.278254710243995e+17, 1.278254710343995e+17, 1.278254710443995e+17, 1.278254710543996e+17, 1.278254710643995e+17, 1.278254710743995e+17, 1.278254710843995e+17, 1.278254710943995e+17, 1.278254711043995e+17, 1.278254711143995e+17, 1.278254711243995e+17, 1.278254711343995e+17, 1.278254711443995e+17, 1.278254711543995e+17, 1.278254711643996e+17, 1.278254711743995e+17, 1.278254711843995e+17, 1.278254711943995e+17, 1.278254712043996e+17, 1.278254712143995e+17, 1.278254712243995e+17, 1.278254712343995e+17, 1.278254712443995e+17, 1.278254712543995e+17, 1.278254712643995e+17, 1.278254712743995e+17, 1.278254712843995e+17, 1.278254712943995e+17, 1.278254713043995e+17, 1.278254713143996e+17, 1.278254713243995e+17, 1.278254713343995e+17, 1.278254713443995e+17, 1.278254713543995e+17, 1.278254713643995e+17, 1.278254713743995e+17, 1.278254713843995e+17, 1.278254713943995e+17, 1.278254714043995e+17, 1.278254714143995e+17, 1.278254714243996e+17, 1.278254714343995e+17, 1.278254714443995e+17, 1.278254714543995e+17, 1.278254714643996e+17, 1.278254714743995e+17, 1.278254714843995e+17, 1.278254714943995e+17, 1.278254715043995e+17, 1.278254715143995e+17, 1.278254715243995e+17, 1.278254715343995e+17, 1.278254715443995e+17, 1.278254715543995e+17, 1.278254715643995e+17, 1.278254715743996e+17, 1.278254715843995e+17, 1.278254715943995e+17, 1.278254716043995e+17, 1.278254716143995e+17, 1.278254716243995e+17, 1.278254716343995e+17, 1.278254716443995e+17, 1.278254716543995e+17, 1.278254716643995e+17, 1.278254716743995e+17, 1.278254716843996e+17, 1.278254716943995e+17, 1.278254717043995e+17, 1.278254717143995e+17, 1.278254717243995e+17, 1.278254717343995e+17, 1.278254717443995e+17, 1.278254717543995e+17, 1.278254717643995e+17, 1.278254717743995e+17, 1.278254717843995e+17, 1.278254717943995e+17, 1.278254718043995e+17, 1.278254718143995e+17, 1.278254718243995e+17, 1.278254718343996e+17, 1.278254718443995e+17, 1.278254718543995e+17, 1.278254718643995e+17, 1.278254718743995e+17, 1.278254718843995e+17, 1.278254718943995e+17, 1.278254719043995e+17, 1.278254719143995e+17, 1.278254719243995e+17, 1.278254719343995e+17, 1.278254719443996e+17, 1.278254719543995e+17, 1.278254719643995e+17, 1.278254719743995e+17, 1.278254719843995e+17, 1.278254719943995e+17, 1.278254720043995e+17, 1.278254720143995e+17, 1.278254720243995e+17, 1.278254720343995e+17, 1.278254720443995e+17, 1.278254720543995e+17, 1.278254720643995e+17, 1.278254720743995e+17, 1.278254720843995e+17, 1.278254720943996e+17, 1.278254721043995e+17, 1.278254721143995e+17, 1.278254721243995e+17, 1.278254721343995e+17, 1.278254721443995e+17, 1.278254721543995e+17, 1.278254721643995e+17, 1.278254721743995e+17, 1.278254721843995e+17, 1.278254721943995e+17, 1.278254722043996e+17, 1.278254722143995e+17, 1.278254722243995e+17, 1.278254722343995e+17, 1.278254722443995e+17, 1.278254722543995e+17, 1.278254722643995e+17, 1.278254722743995e+17, 1.278254722843995e+17, 1.278254722943995e+17, 1.278254723043995e+17, 1.278254723143996e+17, 1.278254723243995e+17, 1.278254723343995e+17, 1.278254723443995e+17, 1.278254723543996e+17, 1.278254723643995e+17, 1.278254723743995e+17, 1.278254723843995e+17, 1.278254723943995e+17, 1.278254724043995e+17, 1.278254724143995e+17, 1.278254724243995e+17, 1.278254724343995e+17, 1.278254724443995e+17, 1.278254724543995e+17, 1.278254724643996e+17, 1.278254724743995e+17, 1.278254724843995e+17, 1.278254724943995e+17, 1.278254725043995e+17, 1.278254725143995e+17, 1.278254725243995e+17, 1.278254725343995e+17, 1.278254725443995e+17, 1.278254725543995e+17, 1.278254725643995e+17, 1.278254725743996e+17, 1.278254725843995e+17, 1.278254725943995e+17, 1.278254726043995e+17, 1.278254726143996e+17, 1.278254726243995e+17, 1.278254726343995e+17, 1.278254726443995e+17, 1.278254726543995e+17, 1.278254726643995e+17, 1.278254726743995e+17, 1.278254726843995e+17, 1.278254726943995e+17, 1.278254727043995e+17, 1.278254727143995e+17, 1.278254727243996e+17, 1.278254727343995e+17, 1.278254727443995e+17, 1.278254727543995e+17, 1.278254727643995e+17, 1.278254727743995e+17, 1.278254727843995e+17, 1.278254727943995e+17, 1.278254728043995e+17, 1.278254728143995e+17, 1.278254728243995e+17, 1.278254728343996e+17, 1.278254728443995e+17, 1.278254728543995e+17, 1.278254728643995e+17, 1.278254728743995e+17, 1.278254728843995e+17, 1.278254728943995e+17, 1.278254729043995e+17, 1.278254729143995e+17, 1.278254729243995e+17, 1.278254729343995e+17, 1.278254729443995e+17, 1.278254729543995e+17, 1.278254729643995e+17, 1.278254729743995e+17, 1.278254729843996e+17, 1.278254729943995e+17, 1.278254730043995e+17, 1.278254730143995e+17, 1.278254730243995e+17, 1.278254730343995e+17, 1.278254730443995e+17, 1.278254730543995e+17, 1.278254730643995e+17, 1.278254730743995e+17, 1.278254730843995e+17, 1.278254730943996e+17, 1.278254731043995e+17, 1.278254731143995e+17, 1.278254731243995e+17, 1.278254731343995e+17, 1.278254731443995e+17, 1.278254731543995e+17, 1.278254731643995e+17, 1.278254731743995e+17, 1.278254731843995e+17, 1.278254731943995e+17, 1.278254732043996e+17, 1.278254732143995e+17, 1.278254732243995e+17, 1.278254732343995e+17, 1.278254732443996e+17, 1.278254732543995e+17, 1.278254732643995e+17, 1.278254732743995e+17, 1.278254732843995e+17, 1.278254732943995e+17, 1.278254733043995e+17, 1.278254733143995e+17, 1.278254733243995e+17, 1.278254733343995e+17, 1.278254733443995e+17, 1.278254733543996e+17, 1.278254733643995e+17, 1.278254733743995e+17, 1.278254733843995e+17, 1.278254733943995e+17, 1.278254734043995e+17, 1.278254734143995e+17, 1.278254734243995e+17, 1.278254734343995e+17, 1.278254734443995e+17, 1.278254734543995e+17, 1.278254734643996e+17, 1.278254734743995e+17, 1.278254734843995e+17, 1.278254734943995e+17, 1.278254735043996e+17, 1.278254735143995e+17, 1.278254735243995e+17, 1.278254735343995e+17, 1.278254735443995e+17, 1.278254735543995e+17, 1.278254735643995e+17, 1.278254735743995e+17, 1.278254735843995e+17, 1.278254735943995e+17, 1.278254736043995e+17, 1.278254736143996e+17, 1.278254736243995e+17, 1.278254736343995e+17, 1.278254736443995e+17, 1.278254736543995e+17, 1.278254736643995e+17, 1.278254736743995e+17, 1.278254736843995e+17, 1.278254736943995e+17, 1.278254737043995e+17, 1.278254737143995e+17, 1.278254737243996e+17, 1.278254737343995e+17, 1.278254737443995e+17, 1.278254737543995e+17, 1.278254737643995e+17, 1.278254737743995e+17, 1.278254737843995e+17, 1.278254737943995e+17, 1.278254738043995e+17, 1.278254738143995e+17, 1.278254738243995e+17, 1.278254738343995e+17, 1.278254738443995e+17, 1.278254738543995e+17, 1.278254738643995e+17, 1.278254738743996e+17, 1.278254738843995e+17, 1.278254738943995e+17, 1.278254739043995e+17, 1.278254739143995e+17, 1.278254739243995e+17, 1.278254739343995e+17, 1.278254739443995e+17, 1.278254739543995e+17, 1.278254739643995e+17, 1.278254739743995e+17, 1.278254739843996e+17, 1.278254739943995e+17, 1.278254740043995e+17, 1.278254740143995e+17, 1.278254740243995e+17, 1.278254740343995e+17, 1.278254740443995e+17, 1.278254740543995e+17, 1.278254740643995e+17, 1.278254740743995e+17, 1.278254740843995e+17, 1.278254740943996e+17, 1.278254741043995e+17, 1.278254741143995e+17, 1.278254741243995e+17, 1.278254741343996e+17, 1.278254741443995e+17, 1.278254741543995e+17, 1.278254741643995e+17, 1.278254741743995e+17, 1.278254741843995e+17, 1.278254741943995e+17, 1.278254742043995e+17, 1.278254742143995e+17, 1.278254742243995e+17, 1.278254742343995e+17, 1.278254742443996e+17, 1.278254742543995e+17, 1.278254742643995e+17, 1.278254742743995e+17, 1.278254742843995e+17, 1.278254742943995e+17, 1.278254743043995e+17, 1.278254743143995e+17, 1.278254743243995e+17, 1.278254743343995e+17, 1.278254743443995e+17, 1.278254743543996e+17, 1.278254743643995e+17, 1.278254743743995e+17, 1.278254743843995e+17, 1.278254743943996e+17, 1.278254744043995e+17, 1.278254744143995e+17, 1.278254744243995e+17, 1.278254744343995e+17, 1.278254744443995e+17, 1.278254744543995e+17, 1.278254744643995e+17, 1.278254744743995e+17, 1.278254744843995e+17, 1.278254744943995e+17, 1.278254745043996e+17, 1.278254745143995e+17, 1.278254745243995e+17, 1.278254745343995e+17, 1.278254745443995e+17, 1.278254745543995e+17, 1.278254745643995e+17, 1.278254745743995e+17, 1.278254745843995e+17, 1.278254745943995e+17, 1.278254746043995e+17, 1.278254746143996e+17, 1.278254746243995e+17, 1.278254746343995e+17, 1.278254746443995e+17, 1.278254746543995e+17, 1.278254746643995e+17, 1.278254746743995e+17, 1.278254746843995e+17, 1.278254746943995e+17, 1.278254747043995e+17, 1.278254747143995e+17, 1.278254747243995e+17, 1.278254747343995e+17, 1.278254747443995e+17, 1.278254747543995e+17, 1.278254747643996e+17, 1.278254747743995e+17, 1.278254747843995e+17, 1.278254747943995e+17, 1.278254748043995e+17, 1.278254748143995e+17, 1.278254748243995e+17, 1.278254748343995e+17, 1.278254748443995e+17, 1.278254748543995e+17, 1.278254748643995e+17, 1.278254748743996e+17, 1.278254748843995e+17, 1.278254748943995e+17, 1.278254749043995e+17, 1.278254749143995e+17, 1.278254749243995e+17, 1.278254749343995e+17, 1.278254749443995e+17, 1.278254749543995e+17, 1.278254749643995e+17, 1.278254749743995e+17, 1.278254749843996e+17, 1.278254749943995e+17, 1.278254750043995e+17, 1.278254750143995e+17, 1.278254750243996e+17, 1.278254750343995e+17, 1.278254750443995e+17, 1.278254750543995e+17, 1.278254750643995e+17, 1.278254750743995e+17, 1.278254750843995e+17, 1.278254750943995e+17, 1.278254751043995e+17, 1.278254751143995e+17, 1.278254751243995e+17, 1.278254751343996e+17, 1.278254751443995e+17, 1.278254751543995e+17, 1.278254751643995e+17, 1.278254751743995e+17, 1.278254751843995e+17, 1.278254751943995e+17, 1.278254752043995e+17, 1.278254752143995e+17, 1.278254752243995e+17, 1.278254752343995e+17, 1.278254752443996e+17, 1.278254752543995e+17, 1.278254752643995e+17, 1.278254752743995e+17, 1.278254752843996e+17, 1.278254752943995e+17, 1.278254753043995e+17, 1.278254753143995e+17, 1.278254753243995e+17, 1.278254753343995e+17, 1.278254753443995e+17, 1.278254753543995e+17, 1.278254753643995e+17, 1.278254753743995e+17, 1.278254753843995e+17, 1.278254753943996e+17, 1.278254754043995e+17, 1.278254754143995e+17, 1.278254754243995e+17, 1.278254754343995e+17, 1.278254754443995e+17, 1.278254754543995e+17, 1.278254754643995e+17, 1.278254754743995e+17, 1.278254754843995e+17, 1.278254754943995e+17, 1.278254755043996e+17, 1.278254755143995e+17, 1.278254755243995e+17, 1.278254755343995e+17, 1.278254755443996e+17, 1.278254755543995e+17, 1.278254755643995e+17, 1.278254755743995e+17, 1.278254755843995e+17, 1.278254755943995e+17, 1.278254756043995e+17, 1.278254756143995e+17, 1.278254756243995e+17, 1.278254756343995e+17, 1.278254756443995e+17, 1.278254756543996e+17, 1.278254756643995e+17, 1.278254756743995e+17, 1.278254756843995e+17, 1.278254756943995e+17, 1.278254757043995e+17, 1.278254757143995e+17, 1.278254757243995e+17, 1.278254757343995e+17, 1.278254757443995e+17, 1.278254757543995e+17, 1.278254757643996e+17, 1.278254757743995e+17, 1.278254757843995e+17, 1.278254757943995e+17, 1.278254758043995e+17, 1.278254758143995e+17, 1.278254758243995e+17, 1.278254758343995e+17, 1.278254758443995e+17, 1.278254758543995e+17, 1.278254758643995e+17, 1.278254758743995e+17, 1.278254758843995e+17, 1.278254758943995e+17, 1.278254759043995e+17, 1.278254759143996e+17, 1.278254759243995e+17, 1.278254759343995e+17, 1.278254759443995e+17, 1.278254759543995e+17, 1.278254759643995e+17, 1.278254759743995e+17, 1.278254759843995e+17, 1.278254759943995e+17, 1.278254760043995e+17, 1.278254760143995e+17, 1.278254760243996e+17, 1.278254760343995e+17, 1.278254760443995e+17, 1.278254760543995e+17, 1.278254760643995e+17, 1.278254760743995e+17, 1.278254760843995e+17, 1.278254760943995e+17, 1.278254761043995e+17, 1.278254761143995e+17, 1.278254761243995e+17, 1.278254761343996e+17, 1.278254761443995e+17, 1.278254761543995e+17, 1.278254761643995e+17, 1.278254761743996e+17, 1.278254761843995e+17, 1.278254761943995e+17, 1.278254762043995e+17, 1.278254762143995e+17, 1.278254762243995e+17, 1.278254762343995e+17, 1.278254762443995e+17, 1.278254762543995e+17, 1.278254762643995e+17, 1.278254762743995e+17, 1.278254762843996e+17, 1.278254762943995e+17, 1.278254763043995e+17, 1.278254763143995e+17, 1.278254763243995e+17, 1.278254763343995e+17, 1.278254763443995e+17, 1.278254763543995e+17, 1.278254763643995e+17, 1.278254763743995e+17, 1.278254763843995e+17, 1.278254763943996e+17, 1.278254764043995e+17, 1.278254764143995e+17, 1.278254764243995e+17, 1.278254764343996e+17, 1.278254764443995e+17, 1.278254764543995e+17, 1.278254764643995e+17, 1.278254764743995e+17, 1.278254764843995e+17, 1.278254764943995e+17, 1.278254765043995e+17, 1.278254765143995e+17, 1.278254765243995e+17, 1.278254765343995e+17, 1.278254765443996e+17, 1.278254765543995e+17, 1.278254765643995e+17, 1.278254765743995e+17, 1.278254765843995e+17, 1.278254765943995e+17, 1.278254766043995e+17, 1.278254766143995e+17, 1.278254766243995e+17, 1.278254766343995e+17, 1.278254766443995e+17, 1.278254766543996e+17, 1.278254766643995e+17, 1.278254766743995e+17, 1.278254766843995e+17, 1.278254766943995e+17, 1.278254767043995e+17, 1.278254767143995e+17, 1.278254767243995e+17, 1.278254767343995e+17, 1.278254767443995e+17, 1.278254767543995e+17, 1.278254767643995e+17, 1.278254767743995e+17, 1.278254767843995e+17, 1.278254767943995e+17, 1.278254768043996e+17, 1.278254768143995e+17, 1.278254768243995e+17, 1.278254768343995e+17, 1.278254768443995e+17, 1.278254768543995e+17, 1.278254768643995e+17, 1.278254768743995e+17, 1.278254768843995e+17, 1.278254768943995e+17, 1.278254769043995e+17, 1.278254769143996e+17, 1.278254769243995e+17, 1.278254769343995e+17, 1.278254769443995e+17, 1.278254769543995e+17, 1.278254769643995e+17, 1.278254769743995e+17, 1.278254769843995e+17, 1.278254769943995e+17, 1.278254770043995e+17, 1.278254770143995e+17, 1.278254770243996e+17, 1.278254770343995e+17, 1.278254770443995e+17, 1.278254770543995e+17, 1.278254770643996e+17, 1.278254770743995e+17, 1.278254770843995e+17, 1.278254770943995e+17, 1.278254771043995e+17, 1.278254771143995e+17, 1.278254771243995e+17, 1.278254771343995e+17, 1.278254771443995e+17, 1.278254771543995e+17, 1.278254771643995e+17, 1.278254771743996e+17, 1.278254771843995e+17, 1.278254771943995e+17, 1.278254772043995e+17, 1.278254772143995e+17, 1.278254772243995e+17, 1.278254772343995e+17, 1.278254772443995e+17, 1.278254772543995e+17, 1.278254772643995e+17, 1.278254772743995e+17, 1.278254772843996e+17, 1.278254772943995e+17, 1.278254773043995e+17, 1.278254773143995e+17, 1.278254773243996e+17, 1.278254773343995e+17, 1.278254773443995e+17, 1.278254773543995e+17, 1.278254773643995e+17, 1.278254773743995e+17, 1.278254773843995e+17, 1.278254773943995e+17, 1.278254774043995e+17, 1.278254774143995e+17, 1.278254774243995e+17, 1.278254774343996e+17, 1.278254774443995e+17, 1.278254774543995e+17, 1.278254774643995e+17, 1.278254774743995e+17, 1.278254774843995e+17, 1.278254774943995e+17, 1.278254775043995e+17, 1.278254775143995e+17, 1.278254775243995e+17, 1.278254775343995e+17, 1.278254775443996e+17, 1.278254775543995e+17, 1.278254775643995e+17, 1.278254775743995e+17, 1.278254775843995e+17, 1.278254775943995e+17, 1.278254776043995e+17, 1.278254776143995e+17, 1.278254776243995e+17, 1.278254776343995e+17, 1.278254776443995e+17, 1.278254776543995e+17, 1.278254776643995e+17, 1.278254776743995e+17, 1.278254776843995e+17, 1.278254776943996e+17, 1.278254777043995e+17, 1.278254777143995e+17, 1.278254777243995e+17, 1.278254777343995e+17, 1.278254777443995e+17, 1.278254777543995e+17, 1.278254777643995e+17, 1.278254777743995e+17, 1.278254777843995e+17, 1.278254777943995e+17, 1.278254778043996e+17, 1.278254778143995e+17, 1.278254778243995e+17, 1.278254778343995e+17, 1.278254778443995e+17, 1.278254778543995e+17, 1.278254778643995e+17, 1.278254778743995e+17, 1.278254778843995e+17, 1.278254778943995e+17, 1.278254779043995e+17, 1.278254779143996e+17, 1.278254779243995e+17, 1.278254779343995e+17, 1.278254779443995e+17, 1.278254779543996e+17, 1.278254779643995e+17, 1.278254779743995e+17, 1.278254779843995e+17, 1.278254779943995e+17, 1.278254780043995e+17, 1.278254780157595e+17, 1.278254780257595e+17, 1.278254780357595e+17, 1.278254780457595e+17, 1.278254780557595e+17, 1.278254780657595e+17, 1.278254780757595e+17, 1.278254780857595e+17, 1.278254780957595e+17, 1.278254781057595e+17, 1.278254781157595e+17, 1.278254781257595e+17, 1.278254781357595e+17, 1.278254781457595e+17, 1.278254781557596e+17, 1.278254781657595e+17, 1.278254781757595e+17, 1.278254781857595e+17, 1.278254781957595e+17, 1.278254782057595e+17, 1.278254782157595e+17, 1.278254782257595e+17, 1.278254782357595e+17, 1.278254782457595e+17, 1.278254782557595e+17, 1.278254782657596e+17, 1.278254782757595e+17, 1.278254782857595e+17, 1.278254782957595e+17, 1.278254783057595e+17, 1.278254783157595e+17, 1.278254783257595e+17, 1.278254783357595e+17, 1.278254783457595e+17, 1.278254783557595e+17, 1.278254783657595e+17, 1.278254783757595e+17, 1.278254783857595e+17, 1.278254783957595e+17, 1.278254784057595e+17, 1.278254784157596e+17, 1.278254784257595e+17, 1.278254784357595e+17, 1.278254784457595e+17, 1.278254784557595e+17, 1.278254784657595e+17, 1.278254784757595e+17, 1.278254784857595e+17, 1.278254784957595e+17, 1.278254785057595e+17, 1.278254785157595e+17, 1.278254785257596e+17, 1.278254785357595e+17, 1.278254785457595e+17, 1.278254785557595e+17, 1.278254785657595e+17, 1.278254785757595e+17, 1.278254785857595e+17, 1.278254785957595e+17, 1.278254786057595e+17, 1.278254786157595e+17, 1.278254786257595e+17, 1.278254786357595e+17, 1.278254786457595e+17, 1.278254786557595e+17, 1.278254786657595e+17, 1.278254786757596e+17, 1.278254786857595e+17, 1.278254786957595e+17, 1.278254787057595e+17, 1.278254787157595e+17, 1.278254787257595e+17, 1.278254787357595e+17, 1.278254787457595e+17, 1.278254787557595e+17, 1.278254787657595e+17, 1.278254787757595e+17, 1.278254787857596e+17, 1.278254787957595e+17, 1.278254788057595e+17, 1.278254788157595e+17, 1.278254788257595e+17, 1.278254788357595e+17, 1.278254788457595e+17, 1.278254788557595e+17, 1.278254788657595e+17, 1.278254788757595e+17, 1.278254788857595e+17, 1.278254788957596e+17, 1.278254789057595e+17, 1.278254789157595e+17, 1.278254789257595e+17, 1.278254789357595e+17, 1.278254789457595e+17, 1.278254789557595e+17, 1.278254789657595e+17, 1.278254789757595e+17, 1.278254789857595e+17, 1.278254789957595e+17, 1.278254790057595e+17, 1.278254790157595e+17, 1.278254790257595e+17, 1.278254790357595e+17, 1.278254790457596e+17, 1.278254790557595e+17, 1.278254790657595e+17, 1.278254790757595e+17, 1.278254790857595e+17, 1.278254790957595e+17, 1.278254791057595e+17, 1.278254791157595e+17, 1.278254791257595e+17, 1.278254791357595e+17, 1.278254791457595e+17, 1.278254791557596e+17, 1.278254791657595e+17, 1.278254791757595e+17, 1.278254791857595e+17, 1.278254791957595e+17, 1.278254792057595e+17, 1.278254792157595e+17, 1.278254792257595e+17, 1.278254792357595e+17, 1.278254792457595e+17, 1.278254792557595e+17, 1.278254792657595e+17, 1.278254792757595e+17, 1.278254792857595e+17, 1.278254792957595e+17, 1.278254793057596e+17, 1.278254793157595e+17, 1.278254793257595e+17, 1.278254793357595e+17, 1.278254793457595e+17, 1.278254793557595e+17, 1.278254793657595e+17, 1.278254793757595e+17, 1.278254793857595e+17, 1.278254793957595e+17, 1.278254794057595e+17, 1.278254794157596e+17, 1.278254794257595e+17, 1.278254794357595e+17, 1.278254794457595e+17, 1.278254794557595e+17, 1.278254794657595e+17, 1.278254794757595e+17, 1.278254794857595e+17, 1.278254794957595e+17, 1.278254795057595e+17, 1.278254795157595e+17, 1.278254795257595e+17, 1.278254795357595e+17, 1.278254795457595e+17, 1.278254795557595e+17, 1.278254795657596e+17, 1.278254795757595e+17, 1.278254795857595e+17, 1.278254795957595e+17, 1.278254796057595e+17, 1.278254796157595e+17, 1.278254796257595e+17, 1.278254796357595e+17, 1.278254796457595e+17, 1.278254796557595e+17, 1.278254796657595e+17, 1.278254796757596e+17, 1.278254796857595e+17, 1.278254796957595e+17, 1.278254797057595e+17, 1.278254797157595e+17, 1.278254797257595e+17, 1.278254797357595e+17, 1.278254797457595e+17, 1.278254797557595e+17, 1.278254797657595e+17, 1.278254797757595e+17, 1.278254797857596e+17, 1.278254797957595e+17, 1.278254798057595e+17, 1.278254798157595e+17, 1.278254798257596e+17, 1.278254798357595e+17, 1.278254798457595e+17, 1.278254798557595e+17, 1.278254798657595e+17, 1.278254798757595e+17, 1.278254798857595e+17, 1.278254798957595e+17, 1.278254799057595e+17, 1.278254799157595e+17, 1.278254799257595e+17, 1.278254799357596e+17, 1.278254799457595e+17, 1.278254799557595e+17, 1.278254799657595e+17, 1.278254799757595e+17, 1.278254799857595e+17, 1.278254799957595e+17, 1.278254800057595e+17, 1.278254800157595e+17, 1.278254800257595e+17, 1.278254800357595e+17, 1.278254800457596e+17, 1.278254800557595e+17, 1.278254800657595e+17, 1.278254800757595e+17, 1.278254800857595e+17, 1.278254800957595e+17, 1.278254801057595e+17, 1.278254801157595e+17, 1.278254801257595e+17, 1.278254801357595e+17, 1.278254801457595e+17, 1.278254801557595e+17, 1.278254801657595e+17, 1.278254801757595e+17, 1.278254801857595e+17, 1.278254801957596e+17, 1.278254802057595e+17, 1.278254802157595e+17, 1.278254802257595e+17, 1.278254802357595e+17, 1.278254802457595e+17, 1.278254802557595e+17, 1.278254802657595e+17, 1.278254802757595e+17, 1.278254802857595e+17, 1.278254802957595e+17, 1.278254803057596e+17, 1.278254803157595e+17, 1.278254803257595e+17, 1.278254803357595e+17, 1.278254803457595e+17, 1.278254803557595e+17, 1.278254803657595e+17, 1.278254803757595e+17, 1.278254803857595e+17, 1.278254803957595e+17, 1.278254804057595e+17, 1.278254804157595e+17, 1.278254804257595e+17, 1.278254804357595e+17, 1.278254804457595e+17, 1.278254804557596e+17, 1.278254804657595e+17, 1.278254804757595e+17, 1.278254804857595e+17, 1.278254804957595e+17, 1.278254805057595e+17, 1.278254805157595e+17, 1.278254805257595e+17, 1.278254805357595e+17, 1.278254805457595e+17, 1.278254805557595e+17, 1.278254805657596e+17, 1.278254805757595e+17, 1.278254805857595e+17, 1.278254805957595e+17, 1.278254806057595e+17, 1.278254806157595e+17, 1.278254806257595e+17, 1.278254806357595e+17, 1.278254806457595e+17, 1.278254806557595e+17, 1.278254806657595e+17, 1.278254806757596e+17, 1.278254806857595e+17, 1.278254806957595e+17, 1.278254807057595e+17, 1.278254807157596e+17, 1.278254807257595e+17, 1.278254807357595e+17, 1.278254807457595e+17, 1.278254807557595e+17, 1.278254807657595e+17, 1.278254807757595e+17, 1.278254807857595e+17, 1.278254807957595e+17, 1.278254808057595e+17, 1.278254808157595e+17, 1.278254808257596e+17, 1.278254808357595e+17, 1.278254808457595e+17, 1.278254808557595e+17, 1.278254808657595e+17, 1.278254808757595e+17, 1.278254808857595e+17, 1.278254808957595e+17, 1.278254809057595e+17, 1.278254809157595e+17, 1.278254809257595e+17, 1.278254809357596e+17, 1.278254809457595e+17, 1.278254809557595e+17, 1.278254809657595e+17, 1.278254809757595e+17, 1.278254809857595e+17, 1.278254809957595e+17, 1.278254810057595e+17, 1.278254810157595e+17, 1.278254810257595e+17, 1.278254810357595e+17, 1.278254810457595e+17, 1.278254810557595e+17, 1.278254810657595e+17, 1.278254810757595e+17, 1.278254810857596e+17, 1.278254810957595e+17, 1.278254811057595e+17, 1.278254811157595e+17, 1.278254811257595e+17, 1.278254811357595e+17, 1.278254811457595e+17, 1.278254811557595e+17, 1.278254811657595e+17, 1.278254811757595e+17, 1.278254811857595e+17, 1.278254811957596e+17, 1.278254812057595e+17, 1.278254812157595e+17, 1.278254812257595e+17, 1.278254812357595e+17, 1.278254812457595e+17, 1.278254812557595e+17, 1.278254812657595e+17, 1.278254812757595e+17, 1.278254812857595e+17, 1.278254812957595e+17, 1.278254813057595e+17, 1.278254813157595e+17, 1.278254813257595e+17, 1.278254813357595e+17, 1.278254813457596e+17, 1.278254813557595e+17, 1.278254813657595e+17, 1.278254813757595e+17, 1.278254813857595e+17, 1.278254813957595e+17, 1.278254814057595e+17, 1.278254814157595e+17, 1.278254814257595e+17, 1.278254814357595e+17, 1.278254814457595e+17, 1.278254814557596e+17, 1.278254814657595e+17, 1.278254814757595e+17, 1.278254814857595e+17, 1.278254814957595e+17, 1.278254815057595e+17, 1.278254815157595e+17, 1.278254815257595e+17, 1.278254815357595e+17, 1.278254815457595e+17, 1.278254815557595e+17, 1.278254815657595e+17, 1.278254815757595e+17, 1.278254815857595e+17, 1.278254815957595e+17, 1.278254816057596e+17, 1.278254816157595e+17, 1.278254816257595e+17, 1.278254816357595e+17, 1.278254816457595e+17, 1.278254816557595e+17, 1.278254816657595e+17, 1.278254816757595e+17, 1.278254816857595e+17, 1.278254816957595e+17, 1.278254817057595e+17, 1.278254817157596e+17, 1.278254817257595e+17, 1.278254817357595e+17, 1.278254817457595e+17, 1.278254817557595e+17, 1.278254817657595e+17, 1.278254817757595e+17, 1.278254817857595e+17, 1.278254817957595e+17, 1.278254818057595e+17, 1.278254818157595e+17, 1.278254818257596e+17, 1.278254818357595e+17, 1.278254818457595e+17, 1.278254818557595e+17, 1.278254818657595e+17, 1.278254818757595e+17, 1.278254818857595e+17, 1.278254818957595e+17, 1.278254819057595e+17, 1.278254819157595e+17, 1.278254819257595e+17, 1.278254819357595e+17, 1.278254819457595e+17, 1.278254819557595e+17, 1.278254819657595e+17, 1.278254819757596e+17, 1.278254819857595e+17, 1.278254819957595e+17, 1.278254820057595e+17, 1.278254820157595e+17, 1.278254820257595e+17, 1.278254820357595e+17, 1.278254820457595e+17, 1.278254820557595e+17, 1.278254820657595e+17, 1.278254820757595e+17, 1.278254820857596e+17, 1.278254820957595e+17, 1.278254821057595e+17, 1.278254821157595e+17, 1.278254821257595e+17, 1.278254821357595e+17, 1.278254821457595e+17, 1.278254821557595e+17, 1.278254821657595e+17, 1.278254821757595e+17, 1.278254821857595e+17, 1.278254821957595e+17, 1.278254822057595e+17, 1.278254822157595e+17, 1.278254822257595e+17, 1.278254822357596e+17, 1.278254822457595e+17, 1.278254822557595e+17, 1.278254822657595e+17, 1.278254822757595e+17, 1.278254822857595e+17, 1.278254822957595e+17, 1.278254823057595e+17, 1.278254823157595e+17, 1.278254823257595e+17, 1.278254823357595e+17, 1.278254823457596e+17, 1.278254823557595e+17, 1.278254823657595e+17, 1.278254823757595e+17, 1.278254823857595e+17, 1.278254823957595e+17, 1.278254824057595e+17, 1.278254824157595e+17, 1.278254824257595e+17, 1.278254824357595e+17, 1.278254824457595e+17, 1.278254824557595e+17, 1.278254824657595e+17, 1.278254824757595e+17, 1.278254824857595e+17, 1.278254824957596e+17, 1.278254825057595e+17, 1.278254825157595e+17, 1.278254825257595e+17, 1.278254825357595e+17, 1.278254825457595e+17, 1.278254825557595e+17, 1.278254825657595e+17, 1.278254825757595e+17, 1.278254825857595e+17, 1.278254825957595e+17, 1.278254826057596e+17, 1.278254826157595e+17, 1.278254826257595e+17, 1.278254826357595e+17, 1.278254826457595e+17, 1.278254826557595e+17, 1.278254826657595e+17, 1.278254826757595e+17, 1.278254826857595e+17, 1.278254826957595e+17, 1.278254827057595e+17, 1.278254827157596e+17, 1.278254827257595e+17, 1.278254827357595e+17, 1.278254827457595e+17, 1.278254827557596e+17, 1.278254827657595e+17, 1.278254827757595e+17, 1.278254827857595e+17, 1.278254827957595e+17, 1.278254828057595e+17, 1.278254828157595e+17, 1.278254828257595e+17, 1.278254828357595e+17, 1.278254828457595e+17, 1.278254828557595e+17, 1.278254828657596e+17, 1.278254828757595e+17, 1.278254828857595e+17, 1.278254828957595e+17, 1.278254829057595e+17, 1.278254829157595e+17, 1.278254829257595e+17, 1.278254829357595e+17, 1.278254829457595e+17, 1.278254829557595e+17, 1.278254829657595e+17, 1.278254829757596e+17, 1.278254829857595e+17, 1.278254829957595e+17, 1.278254830057595e+17, 1.278254830157595e+17, 1.278254830257595e+17, 1.278254830357595e+17, 1.278254830457595e+17, 1.278254830557595e+17, 1.278254830657595e+17, 1.278254830757595e+17, 1.278254830857595e+17, 1.278254830957595e+17, 1.278254831057595e+17, 1.278254831157595e+17, 1.278254831257596e+17, 1.278254831357595e+17, 1.278254831457595e+17, 1.278254831557595e+17, 1.278254831657595e+17, 1.278254831757595e+17, 1.278254831857595e+17, 1.278254831957595e+17, 1.278254832057595e+17, 1.278254832157595e+17, 1.278254832257595e+17, 1.278254832357596e+17, 1.278254832457595e+17, 1.278254832557595e+17, 1.278254832657595e+17, 1.278254832757595e+17, 1.278254832857595e+17, 1.278254832957595e+17, 1.278254833057595e+17, 1.278254833157595e+17, 1.278254833257595e+17, 1.278254833357595e+17, 1.278254833457595e+17, 1.278254833557595e+17, 1.278254833657595e+17, 1.278254833757595e+17, 1.278254833857596e+17, 1.278254833957595e+17, 1.278254834057595e+17, 1.278254834157595e+17, 1.278254834257595e+17, 1.278254834357595e+17, 1.278254834457595e+17, 1.278254834557595e+17, 1.278254834657595e+17, 1.278254834757595e+17, 1.278254834857595e+17, 1.278254834957596e+17, 1.278254835057595e+17, 1.278254835157595e+17, 1.278254835257595e+17, 1.278254835357595e+17, 1.278254835457595e+17, 1.278254835557595e+17, 1.278254835657595e+17, 1.278254835757595e+17, 1.278254835857595e+17, 1.278254835957595e+17, 1.278254836057596e+17, 1.278254836157595e+17, 1.278254836257595e+17, 1.278254836357595e+17, 1.278254836457596e+17, 1.278254836557595e+17, 1.278254836657595e+17, 1.278254836757595e+17, 1.278254836857595e+17, 1.278254836957595e+17, 1.278254837057595e+17, 1.278254837157595e+17, 1.278254837257595e+17, 1.278254837357595e+17, 1.278254837457595e+17, 1.278254837557596e+17, 1.278254837657595e+17, 1.278254837757595e+17, 1.278254837857595e+17, 1.278254837957595e+17, 1.278254838057595e+17, 1.278254838157595e+17, 1.278254838257595e+17, 1.278254838357595e+17, 1.278254838457595e+17, 1.278254838557595e+17, 1.278254838657596e+17, 1.278254838757595e+17, 1.278254838857595e+17, 1.278254838957595e+17, 1.278254839057595e+17, 1.278254839157595e+17, 1.278254839257595e+17, 1.278254839357595e+17, 1.278254839457595e+17, 1.278254839557595e+17, 1.278254839657595e+17, 1.278254839757595e+17, 1.278254839857595e+17, 1.278254839957595e+17, 1.278254840057595e+17, 1.278254840157596e+17, 1.278254840257595e+17, 1.278254840357595e+17, 1.278254840457595e+17, 1.278254840557595e+17, 1.278254840657595e+17, 1.278254840757595e+17, 1.278254840857595e+17, 1.278254840957595e+17, 1.278254841057595e+17, 1.278254841157595e+17, 1.278254841257596e+17, 1.278254841357595e+17, 1.278254841457595e+17, 1.278254841557595e+17, 1.278254841657595e+17, 1.278254841757595e+17, 1.278254841857595e+17, 1.278254841957595e+17, 1.278254842057595e+17, 1.278254842157595e+17, 1.278254842257595e+17, 1.278254842357595e+17, 1.278254842457595e+17, 1.278254842557595e+17, 1.278254842657595e+17, 1.278254842757596e+17, 1.278254842857595e+17, 1.278254842957595e+17, 1.278254843057595e+17, 1.278254843157595e+17, 1.278254843257595e+17, 1.278254843357595e+17, 1.278254843457595e+17, 1.278254843557595e+17, 1.278254843657595e+17, 1.278254843757595e+17, 1.278254843857596e+17, 1.278254843957595e+17, 1.278254844057595e+17, 1.278254844157595e+17, 1.278254844257595e+17, 1.278254844357595e+17, 1.278254844457595e+17, 1.278254844557595e+17, 1.278254844657595e+17, 1.278254844757595e+17, 1.278254844857595e+17, 1.278254844957595e+17, 1.278254845057595e+17, 1.278254845157595e+17, 1.278254845257595e+17, 1.278254845357596e+17, 1.278254845457595e+17, 1.278254845557595e+17, 1.278254845657595e+17, 1.278254845757595e+17, 1.278254845857595e+17, 1.278254845957595e+17, 1.278254846057595e+17, 1.278254846157595e+17, 1.278254846257595e+17, 1.278254846357595e+17, 1.278254846457596e+17, 1.278254846557595e+17, 1.278254846657595e+17, 1.278254846757595e+17, 1.278254846857595e+17, 1.278254846957595e+17, 1.278254847057595e+17, 1.278254847157595e+17, 1.278254847257595e+17, 1.278254847357595e+17, 1.278254847457595e+17, 1.278254847557596e+17, 1.278254847657595e+17, 1.278254847757595e+17, 1.278254847857595e+17, 1.278254847957595e+17, 1.278254848057595e+17, 1.278254848157595e+17, 1.278254848257595e+17, 1.278254848357595e+17, 1.278254848457595e+17, 1.278254848557595e+17, 1.278254848657595e+17, 1.278254848757595e+17, 1.278254848857595e+17, 1.278254848957595e+17, 1.278254849057596e+17, 1.278254849157595e+17, 1.278254849257595e+17, 1.278254849357595e+17, 1.278254849457595e+17, 1.278254849557595e+17, 1.278254849657595e+17, 1.278254849757595e+17, 1.278254849857595e+17, 1.278254849957595e+17, 1.278254850057595e+17, 1.278254850157596e+17, 1.278254850257595e+17, 1.278254850357595e+17, 1.278254850457595e+17, 1.278254850557595e+17, 1.278254850657595e+17, 1.278254850757595e+17, 1.278254850857595e+17, 1.278254850957595e+17, 1.278254851057595e+17, 1.278254851157595e+17, 1.278254851257595e+17, 1.278254851357595e+17, 1.278254851457595e+17, 1.278254851557595e+17, 1.278254851657596e+17, 1.278254851757595e+17, 1.278254851857595e+17, 1.278254851957595e+17, 1.278254852057595e+17, 1.278254852157595e+17, 1.278254852257595e+17, 1.278254852357595e+17, 1.278254852457595e+17, 1.278254852557595e+17, 1.278254852657595e+17, 1.278254852757596e+17, 1.278254852857595e+17, 1.278254852957595e+17, 1.278254853057595e+17, 1.278254853157595e+17, 1.278254853257595e+17, 1.278254853357595e+17, 1.278254853457595e+17, 1.278254853557595e+17, 1.278254853657595e+17, 1.278254853757595e+17, 1.278254853857595e+17, 1.278254853957595e+17, 1.278254854057595e+17, 1.278254854157595e+17, 1.278254854257596e+17, 1.278254854357595e+17, 1.278254854457595e+17, 1.278254854557595e+17, 1.278254854657595e+17, 1.278254854757595e+17, 1.278254854857595e+17, 1.278254854957595e+17, 1.278254855057595e+17, 1.278254855157595e+17, 1.278254855257595e+17, 1.278254855357596e+17, 1.278254855457595e+17, 1.278254855557595e+17, 1.278254855657595e+17, 1.278254855757595e+17, 1.278254855857595e+17, 1.278254855957595e+17, 1.278254856057595e+17, 1.278254856157595e+17, 1.278254856257595e+17, 1.278254856357595e+17, 1.278254856457596e+17, 1.278254856557595e+17, 1.278254856657595e+17, 1.278254856757595e+17, 1.278254856857595e+17, 1.278254856957595e+17, 1.278254857057595e+17, 1.278254857157595e+17, 1.278254857257595e+17, 1.278254857357595e+17, 1.278254857457595e+17, 1.278254857557595e+17, 1.278254857657595e+17, 1.278254857757595e+17, 1.278254857857595e+17, 1.278254857957596e+17, 1.278254858057595e+17, 1.278254858157595e+17, 1.278254858257595e+17, 1.278254858357595e+17, 1.278254858457595e+17, 1.278254858557595e+17, 1.278254858657595e+17, 1.278254858757595e+17, 1.278254858857595e+17, 1.278254858957595e+17, 1.278254859057596e+17, 1.278254859157595e+17, 1.278254859257595e+17, 1.278254859357595e+17, 1.278254859457595e+17, 1.278254859557595e+17, 1.278254859657595e+17, 1.278254859757595e+17, 1.278254859857595e+17, 1.278254859957595e+17, 1.278254860057595e+17, 1.278254860157595e+17, 1.278254860257595e+17, 1.278254860357595e+17, 1.278254860457595e+17, 1.278254860557596e+17, 1.278254860657595e+17, 1.278254860757595e+17, 1.278254860857595e+17, 1.278254860957595e+17, 1.278254861057595e+17, 1.278254861157595e+17, 1.278254861257595e+17, 1.278254861357595e+17, 1.278254861457595e+17, 1.278254861557595e+17, 1.278254861657596e+17, 1.278254861757595e+17, 1.278254861857595e+17, 1.278254861957595e+17, 1.278254862057595e+17, 1.278254862157595e+17, 1.278254862257595e+17, 1.278254862357595e+17, 1.278254862457595e+17, 1.278254862557595e+17, 1.278254862657595e+17, 1.278254862757595e+17, 1.278254862857595e+17, 1.278254862957595e+17, 1.278254863057595e+17, 1.278254863157596e+17, 1.278254863257595e+17, 1.278254863357595e+17, 1.278254863457595e+17, 1.278254863557595e+17, 1.278254863657595e+17, 1.278254863757595e+17, 1.278254863857595e+17, 1.278254863957595e+17, 1.278254864057595e+17, 1.278254864157595e+17, 1.278254864257596e+17, 1.278254864357595e+17, 1.278254864457595e+17, 1.278254864557595e+17, 1.278254864657595e+17, 1.278254864757595e+17, 1.278254864857595e+17, 1.278254864957595e+17, 1.278254865057595e+17, 1.278254865157595e+17, 1.278254865257595e+17, 1.278254865357596e+17, 1.278254865457595e+17, 1.278254865557595e+17, 1.278254865657595e+17, 1.278254865757596e+17, 1.278254865857595e+17, 1.278254865957595e+17, 1.278254866057595e+17, 1.278254866157595e+17, 1.278254866257595e+17, 1.278254866357595e+17, 1.278254866457595e+17, 1.278254866557595e+17, 1.278254866657595e+17, 1.278254866757595e+17, 1.278254866857596e+17, 1.278254866957595e+17, 1.278254867057595e+17, 1.278254867157595e+17, 1.278254867257595e+17, 1.278254867357595e+17, 1.278254867457595e+17, 1.278254867557595e+17, 1.278254867657595e+17, 1.278254867757595e+17, 1.278254867857595e+17, 1.278254867957596e+17, 1.278254868057595e+17, 1.278254868157595e+17, 1.278254868257595e+17, 1.278254868357595e+17, 1.278254868457595e+17, 1.278254868557595e+17, 1.278254868657595e+17, 1.278254868757595e+17, 1.278254868857595e+17, 1.278254868957595e+17, 1.278254869057595e+17, 1.278254869157595e+17, 1.278254869257595e+17, 1.278254869357595e+17, 1.278254869457596e+17, 1.278254869557595e+17, 1.278254869657595e+17, 1.278254869757595e+17, 1.278254869857595e+17, 1.278254869957595e+17, 1.278254870057595e+17, 1.278254870157595e+17, 1.278254870257595e+17, 1.278254870357595e+17, 1.278254870457595e+17, 1.278254870557596e+17, 1.278254870657595e+17, 1.278254870757595e+17, 1.278254870857595e+17, 1.278254870957595e+17, 1.278254871057595e+17, 1.278254871157595e+17, 1.278254871257595e+17, 1.278254871357595e+17, 1.278254871457595e+17, 1.278254871557595e+17, 1.278254871657595e+17, 1.278254871757595e+17, 1.278254871857595e+17, 1.278254871957595e+17, 1.278254872057596e+17, 1.278254872157595e+17, 1.278254872257595e+17, 1.278254872357595e+17, 1.278254872457595e+17, 1.278254872557595e+17, 1.278254872657595e+17, 1.278254872757595e+17, 1.278254872857595e+17, 1.278254872957595e+17, 1.278254873057595e+17, 1.278254873157596e+17, 1.278254873257595e+17, 1.278254873357595e+17, 1.278254873457595e+17, 1.278254873557595e+17, 1.278254873657595e+17, 1.278254873757595e+17, 1.278254873857595e+17, 1.278254873957595e+17, 1.278254874057595e+17, 1.278254874157595e+17, 1.278254874257596e+17, 1.278254874357595e+17, 1.278254874457595e+17, 1.278254874557595e+17, 1.278254874657596e+17, 1.278254874757595e+17, 1.278254874857595e+17, 1.278254874957595e+17, 1.278254875057595e+17, 1.278254875157595e+17, 1.278254875257595e+17, 1.278254875357595e+17, 1.278254875457595e+17, 1.278254875557595e+17, 1.278254875657595e+17, 1.278254875757596e+17, 1.278254875857595e+17, 1.278254875957595e+17, 1.278254876057595e+17, 1.278254876157595e+17, 1.278254876257595e+17, 1.278254876357595e+17, 1.278254876457595e+17, 1.278254876557595e+17, 1.278254876657595e+17, 1.278254876757595e+17, 1.278254876857596e+17, 1.278254876957595e+17, 1.278254877057595e+17, 1.278254877157595e+17, 1.278254877257595e+17, 1.278254877357595e+17, 1.278254877457595e+17, 1.278254877557595e+17, 1.278254877657595e+17, 1.278254877757595e+17, 1.278254877857595e+17, 1.278254877957595e+17, 1.278254878057595e+17, 1.278254878157595e+17, 1.278254878257595e+17, 1.278254878357596e+17, 1.278254878457595e+17, 1.278254878557595e+17, 1.278254878657595e+17, 1.278254878757595e+17, 1.278254878857595e+17, 1.278254878957595e+17, 1.278254879057595e+17, 1.278254879157595e+17, 1.278254879257595e+17, 1.278254879357595e+17, 1.278254879457596e+17, 1.278254879557595e+17, 1.278254879657595e+17, 1.278254879757595e+17, 1.278254879857595e+17, 1.278254879957595e+17, 1.278254880057595e+17, 1.278254880157595e+17, 1.278254880257595e+17, 1.278254880357595e+17, 1.278254880457595e+17, 1.278254880557595e+17, 1.278254880657595e+17, 1.278254880757595e+17, 1.278254880857595e+17, 1.278254880957596e+17, 1.278254881057595e+17, 1.278254881157595e+17, 1.278254881257595e+17, 1.278254881357595e+17, 1.278254881457595e+17, 1.278254881557595e+17, 1.278254881657595e+17, 1.278254881757595e+17, 1.278254881857595e+17, 1.278254881957595e+17, 1.278254882057596e+17, 1.278254882157595e+17, 1.278254882257595e+17, 1.278254882357595e+17, 1.278254882457595e+17, 1.278254882557595e+17, 1.278254882657595e+17, 1.278254882757595e+17, 1.278254882857595e+17, 1.278254882957595e+17, 1.278254883057595e+17, 1.278254883157595e+17, 1.278254883257595e+17, 1.278254883357595e+17, 1.278254883457595e+17, 1.278254883557596e+17, 1.278254883657595e+17, 1.278254883757595e+17, 1.278254883857595e+17, 1.278254883957595e+17, 1.278254884057595e+17, 1.278254884157595e+17, 1.278254884257595e+17, 1.278254884357595e+17, 1.278254884457595e+17, 1.278254884557595e+17, 1.278254884657596e+17, 1.278254884757595e+17, 1.278254884857595e+17, 1.278254884957595e+17, 1.278254885057595e+17, 1.278254885157595e+17, 1.278254885257595e+17, 1.278254885357595e+17, 1.278254885457595e+17, 1.278254885557595e+17, 1.278254885657595e+17, 1.278254885757596e+17, 1.278254885857595e+17, 1.278254885957595e+17, 1.278254886057595e+17, 1.278254886157595e+17, 1.278254886257595e+17, 1.278254886357595e+17, 1.278254886457595e+17, 1.278254886557595e+17, 1.278254886657595e+17, 1.278254886757595e+17, 1.278254886857595e+17, 1.278254886957595e+17, 1.278254887057595e+17, 1.278254887157595e+17, 1.278254887257596e+17, 1.278254887357595e+17, 1.278254887457595e+17, 1.278254887557595e+17, 1.278254887657595e+17, 1.278254887757595e+17, 1.278254887857595e+17, 1.278254887957595e+17, 1.278254888057595e+17, 1.278254888157595e+17, 1.278254888257595e+17, 1.278254888357596e+17, 1.278254888457595e+17, 1.278254888557595e+17, 1.278254888657595e+17, 1.278254888757595e+17, 1.278254888857595e+17, 1.278254888957595e+17, 1.278254889057595e+17, 1.278254889157595e+17, 1.278254889257595e+17, 1.278254889357595e+17, 1.278254889457595e+17, 1.278254889557595e+17, 1.278254889657595e+17, 1.278254889757595e+17, 1.278254889857596e+17, 1.278254889957595e+17, 1.278254890057595e+17, 1.278254890157595e+17, 1.278254890257595e+17, 1.278254890357595e+17, 1.278254890457595e+17, 1.278254890557595e+17, 1.278254890657595e+17, 1.278254890757595e+17, 1.278254890857595e+17, 1.278254890957596e+17, 1.278254891057595e+17, 1.278254891157595e+17, 1.278254891257595e+17, 1.278254891357595e+17, 1.278254891457595e+17, 1.278254891557595e+17, 1.278254891657595e+17, 1.278254891757595e+17, 1.278254891857595e+17, 1.278254891957595e+17, 1.278254892057595e+17, 1.278254892157595e+17, 1.278254892257595e+17, 1.278254892357595e+17, 1.278254892457596e+17, 1.278254892557595e+17, 1.278254892657595e+17, 1.278254892757595e+17, 1.278254892857595e+17, 1.278254892957595e+17, 1.278254893057595e+17, 1.278254893157595e+17, 1.278254893257595e+17, 1.278254893357595e+17, 1.278254893457595e+17, 1.278254893557596e+17, 1.278254893657595e+17, 1.278254893757595e+17, 1.278254893857595e+17, 1.278254893957595e+17, 1.278254894057595e+17, 1.278254894157595e+17, 1.278254894257595e+17, 1.278254894357595e+17, 1.278254894457595e+17, 1.278254894557595e+17, 1.278254894657596e+17, 1.278254894757595e+17, 1.278254894857595e+17, 1.278254894957595e+17, 1.278254895057596e+17, 1.278254895157595e+17, 1.278254895257595e+17, 1.278254895357595e+17, 1.278254895457595e+17, 1.278254895557595e+17, 1.278254895657595e+17, 1.278254895757595e+17, 1.278254895857595e+17, 1.278254895957595e+17, 1.278254896057595e+17, 1.278254896157596e+17, 1.278254896257595e+17, 1.278254896357595e+17, 1.278254896457595e+17, 1.278254896557595e+17, 1.278254896657595e+17, 1.278254896757595e+17, 1.278254896857595e+17, 1.278254896957595e+17, 1.278254897057595e+17, 1.278254897157595e+17, 1.278254897257596e+17, 1.278254897357595e+17, 1.278254897457595e+17, 1.278254897557595e+17, 1.278254897657595e+17, 1.278254897757595e+17, 1.278254897857595e+17, 1.278254897957595e+17, 1.278254898057595e+17, 1.278254898157595e+17, 1.278254898257595e+17, 1.278254898357595e+17, 1.278254898457595e+17, 1.278254898557595e+17, 1.278254898657595e+17, 1.278254898757596e+17, 1.278254898857595e+17, 1.278254898957595e+17, 1.278254899057595e+17, 1.278254899157595e+17, 1.278254899257595e+17, 1.278254899357595e+17, 1.278254899457595e+17, 1.278254899557595e+17, 1.278254899657595e+17, 1.278254899757595e+17, 1.278254899857596e+17, 1.278254899957595e+17, 1.278254900057595e+17, 1.278254900157595e+17, 1.278254900257595e+17, 1.278254900357595e+17, 1.278254900457595e+17, 1.278254900557595e+17, 1.278254900657595e+17, 1.278254900757595e+17, 1.278254900857595e+17, 1.278254900957595e+17, 1.278254901057595e+17, 1.278254901157595e+17, 1.278254901257595e+17, 1.278254901357596e+17, 1.278254901457595e+17, 1.278254901557595e+17, 1.278254901657595e+17, 1.278254901757595e+17, 1.278254901857595e+17, 1.278254901957595e+17, 1.278254902057595e+17, 1.278254902157595e+17, 1.278254902257595e+17, 1.278254902357595e+17, 1.278254902457596e+17, 1.278254902557595e+17, 1.278254902657595e+17, 1.278254902757595e+17, 1.278254902857595e+17, 1.278254902957595e+17, 1.278254903057595e+17, 1.278254903157595e+17, 1.278254903257595e+17, 1.278254903357595e+17, 1.278254903457595e+17, 1.278254903557596e+17, 1.278254903657595e+17, 1.278254903757595e+17, 1.278254903857595e+17, 1.278254903957596e+17, 1.278254904057595e+17, 1.278254904157595e+17, 1.278254904257595e+17, 1.278254904357595e+17, 1.278254904457595e+17, 1.278254904557595e+17, 1.278254904657595e+17, 1.278254904757595e+17, 1.278254904857595e+17, 1.278254904957595e+17, 1.278254905057596e+17, 1.278254905157595e+17, 1.278254905257595e+17, 1.278254905357595e+17, 1.278254905457595e+17, 1.278254905557595e+17, 1.278254905657595e+17, 1.278254905757595e+17, 1.278254905857595e+17, 1.278254905957595e+17, 1.278254906057595e+17, 1.278254906157596e+17, 1.278254906257595e+17, 1.278254906357595e+17, 1.278254906457595e+17, 1.278254906557595e+17, 1.278254906657595e+17, 1.278254906757595e+17, 1.278254906857595e+17, 1.278254906957595e+17, 1.278254907057595e+17, 1.278254907157595e+17, 1.278254907257595e+17, 1.278254907357595e+17, 1.278254907457595e+17, 1.278254907557595e+17, 1.278254907657596e+17, 1.278254907757595e+17, 1.278254907857595e+17, 1.278254907957595e+17, 1.278254908057595e+17, 1.278254908157595e+17, 1.278254908257595e+17, 1.278254908357595e+17, 1.278254908457595e+17, 1.278254908557595e+17, 1.278254908657595e+17, 1.278254908757596e+17, 1.278254908857595e+17, 1.278254908957595e+17, 1.278254909057595e+17, 1.278254909157595e+17, 1.278254909257595e+17, 1.278254909357595e+17, 1.278254909457595e+17, 1.278254909557595e+17, 1.278254909657595e+17, 1.278254909757595e+17, 1.278254909857595e+17, 1.278254909957595e+17, 1.278254910057595e+17, 1.278254910157595e+17, 1.278254910257596e+17, 1.278254910357595e+17, 1.278254910457595e+17, 1.278254910557595e+17, 1.278254910657595e+17, 1.278254910757595e+17, 1.278254910857595e+17, 1.278254910957595e+17, 1.278254911057595e+17, 1.278254911157595e+17, 1.278254911257595e+17, 1.278254911357596e+17, 1.278254911457595e+17, 1.278254911557595e+17, 1.278254911657595e+17, 1.278254911757595e+17, 1.278254911857595e+17, 1.278254911957595e+17, 1.278254912057595e+17, 1.278254912157595e+17, 1.278254912257595e+17, 1.278254912357595e+17, 1.278254912457595e+17, 1.278254912557595e+17, 1.278254912657595e+17, 1.278254912757595e+17, 1.278254912857596e+17, 1.278254912957595e+17, 1.278254913057595e+17, 1.278254913157595e+17, 1.278254913257595e+17, 1.278254913357595e+17, 1.278254913457595e+17, 1.278254913557595e+17, 1.278254913657595e+17, 1.278254913757595e+17, 1.278254913857595e+17, 1.278254913957596e+17, 1.278254914057595e+17, 1.278254914157595e+17, 1.278254914257595e+17, 1.278254914357595e+17, 1.278254914457595e+17, 1.278254914557595e+17, 1.278254914657595e+17, 1.278254914757595e+17, 1.278254914857595e+17, 1.278254914957595e+17, 1.278254915057596e+17, 1.278254915157595e+17, 1.278254915257595e+17, 1.278254915357595e+17, 1.278254915457595e+17, 1.278254915557595e+17, 1.278254915657595e+17, 1.278254915757595e+17, 1.278254915857595e+17, 1.278254915957595e+17, 1.278254916057595e+17, 1.278254916157595e+17, 1.278254916257595e+17, 1.278254916357595e+17, 1.278254916457595e+17, 1.278254916557596e+17, 1.278254916657595e+17, 1.278254916757595e+17, 1.278254916857595e+17, 1.278254916957595e+17, 1.278254917057595e+17, 1.278254917157595e+17, 1.278254917257595e+17, 1.278254917357595e+17, 1.278254917457595e+17, 1.278254917557595e+17, 1.278254917657596e+17, 1.278254917757595e+17, 1.278254917857595e+17, 1.278254917957595e+17, 1.278254918057595e+17, 1.278254918157595e+17, 1.278254918257595e+17, 1.278254918357595e+17, 1.278254918457595e+17, 1.278254918557595e+17, 1.278254918657595e+17, 1.278254918757595e+17, 1.278254918857595e+17, 1.278254918957595e+17, 1.278254919057595e+17, 1.278254919157596e+17, 1.278254919257595e+17, 1.278254919357595e+17, 1.278254919457595e+17, 1.278254919557595e+17, 1.278254919657595e+17, 1.278254919757595e+17, 1.278254919857595e+17, 1.278254919957595e+17, 1.278254920057595e+17, 1.278254920157595e+17, 1.278254920257596e+17, 1.278254920357595e+17, 1.278254920457595e+17, 1.278254920557595e+17, 1.278254920657595e+17, 1.278254920757595e+17, 1.278254920857595e+17, 1.278254920957595e+17, 1.278254921057595e+17, 1.278254921157595e+17, 1.278254921257595e+17, 1.278254921357595e+17, 1.278254921457595e+17, 1.278254921557595e+17, 1.278254921657595e+17, 1.278254921757596e+17, 1.278254921857595e+17, 1.278254921957595e+17, 1.278254922057595e+17, 1.278254922157595e+17, 1.278254922257595e+17, 1.278254922357595e+17, 1.278254922457595e+17, 1.278254922557595e+17, 1.278254922657595e+17, 1.278254922757595e+17, 1.278254922857596e+17, 1.278254922957595e+17, 1.278254923057595e+17, 1.278254923157595e+17, 1.278254923257595e+17, 1.278254923357595e+17, 1.278254923457595e+17, 1.278254923557595e+17, 1.278254923657595e+17, 1.278254923757595e+17, 1.278254923857595e+17, 1.278254923957596e+17, 1.278254924057595e+17, 1.278254924157595e+17, 1.278254924257595e+17, 1.278254924357595e+17, 1.278254924457595e+17, 1.278254924557595e+17, 1.278254924657595e+17, 1.278254924757595e+17, 1.278254924857595e+17, 1.278254924957595e+17, 1.278254925057595e+17, 1.278254925157595e+17, 1.278254925257595e+17, 1.278254925357595e+17, 1.278254925457596e+17, 1.278254925557595e+17, 1.278254925657595e+17, 1.278254925757595e+17, 1.278254925857595e+17, 1.278254925957595e+17, 1.278254926057595e+17, 1.278254926157595e+17, 1.278254926257595e+17, 1.278254926357595e+17, 1.278254926457595e+17, 1.278254926557596e+17, 1.278254926657595e+17, 1.278254926757595e+17, 1.278254926857595e+17, 1.278254926957595e+17, 1.278254927057595e+17, 1.278254927157595e+17, 1.278254927257595e+17, 1.278254927357595e+17, 1.278254927457595e+17, 1.278254927557595e+17, 1.278254927657595e+17, 1.278254927757595e+17, 1.278254927857595e+17, 1.278254927957595e+17, 1.278254928057596e+17, 1.278254928157595e+17, 1.278254928257595e+17, 1.278254928357595e+17, 1.278254928457595e+17, 1.278254928557595e+17, 1.278254928657595e+17, 1.278254928757595e+17, 1.278254928857595e+17, 1.278254928957595e+17, 1.278254929057595e+17, 1.278254929157596e+17, 1.278254929257595e+17, 1.278254929357595e+17, 1.278254929457595e+17, 1.278254929557595e+17, 1.278254929657595e+17, 1.278254929757595e+17, 1.278254929857595e+17, 1.278254929957595e+17, 1.278254930057595e+17, 1.278254930157595e+17, 1.278254930257595e+17, 1.278254930357595e+17, 1.278254930457595e+17, 1.278254930557595e+17, 1.278254930657596e+17, 1.278254930757595e+17, 1.278254930857595e+17, 1.278254930957595e+17, 1.278254931057595e+17, 1.278254931157595e+17, 1.278254931257595e+17, 1.278254931357595e+17, 1.278254931457595e+17, 1.278254931557595e+17, 1.278254931657595e+17, 1.278254931757596e+17, 1.278254931857595e+17, 1.278254931957595e+17, 1.278254932057595e+17, 1.278254932157595e+17, 1.278254932257595e+17, 1.278254932357595e+17, 1.278254932457595e+17, 1.278254932557595e+17, 1.278254932657595e+17, 1.278254932757595e+17, 1.278254932857596e+17, 1.278254932957595e+17, 1.278254933057595e+17, 1.278254933157595e+17, 1.278254933257596e+17, 1.278254933357595e+17, 1.278254933457595e+17, 1.278254933557595e+17, 1.278254933657595e+17, 1.278254933757595e+17, 1.278254933857595e+17, 1.278254933957595e+17, 1.278254934057595e+17, 1.278254934157595e+17, 1.278254934257595e+17, 1.278254934357596e+17, 1.278254934457595e+17, 1.278254934557595e+17, 1.278254934657595e+17, 1.278254934757595e+17, 1.278254934857595e+17, 1.278254934957595e+17, 1.278254935057595e+17, 1.278254935157595e+17, 1.278254935257595e+17, 1.278254935357595e+17, 1.278254935457596e+17, 1.278254935557595e+17, 1.278254935657595e+17, 1.278254935757595e+17, 1.278254935857595e+17, 1.278254935957595e+17, 1.278254936057595e+17, 1.278254936157595e+17, 1.278254936257595e+17, 1.278254936357595e+17, 1.278254936457595e+17, 1.278254936557595e+17, 1.278254936657595e+17, 1.278254936757595e+17, 1.278254936857595e+17, 1.278254936957596e+17, 1.278254937057595e+17, 1.278254937157595e+17, 1.278254937257595e+17, 1.278254937357595e+17, 1.278254937457595e+17, 1.278254937557595e+17, 1.278254937657595e+17, 1.278254937757595e+17, 1.278254937857595e+17, 1.278254937957595e+17, 1.278254938057596e+17, 1.278254938157595e+17, 1.278254938257595e+17, 1.278254938357595e+17, 1.278254938457595e+17, 1.278254938557595e+17, 1.278254938657595e+17, 1.278254938757595e+17, 1.278254938857595e+17, 1.278254938957595e+17, 1.278254939057595e+17, 1.278254939157595e+17, 1.278254939257595e+17, 1.278254939357595e+17, 1.278254939457595e+17, 1.278254939557596e+17, 1.278254939657595e+17, 1.278254939757595e+17, 1.278254939857595e+17, 1.278254939957595e+17, 1.278254940057595e+17, 1.278254940157595e+17, 1.278254940257595e+17, 1.278254940357595e+17, 1.278254940457595e+17, 1.278254940557595e+17, 1.278254940657596e+17, 1.278254940757595e+17, 1.278254940857595e+17, 1.278254940957595e+17, 1.278254941057595e+17, 1.278254941157595e+17, 1.278254941257595e+17, 1.278254941357595e+17, 1.278254941457595e+17, 1.278254941557595e+17, 1.278254941657595e+17, 1.278254941757596e+17, 1.278254941857595e+17, 1.278254941957595e+17, 1.278254942057595e+17, 1.278254942157596e+17, 1.278254942257595e+17, 1.278254942357595e+17, 1.278254942457595e+17, 1.278254942557595e+17, 1.278254942657595e+17, 1.278254942757595e+17, 1.278254942857595e+17, 1.278254942957595e+17, 1.278254943057595e+17, 1.278254943157595e+17, 1.278254943257596e+17, 1.278254943357595e+17, 1.278254943457595e+17, 1.278254943557595e+17, 1.278254943657595e+17, 1.278254943757595e+17, 1.278254943857595e+17, 1.278254943957595e+17, 1.278254944057595e+17, 1.278254944157595e+17, 1.278254944257595e+17, 1.278254944357596e+17, 1.278254944457595e+17, 1.278254944557595e+17, 1.278254944657595e+17, 1.278254944757595e+17, 1.278254944857595e+17, 1.278254944957595e+17, 1.278254945057595e+17, 1.278254945157595e+17, 1.278254945257595e+17, 1.278254945357595e+17, 1.278254945457595e+17, 1.278254945557595e+17, 1.278254945657595e+17, 1.278254945757595e+17, 1.278254945857596e+17, 1.278254945957595e+17, 1.278254946057595e+17, 1.278254946157595e+17, 1.278254946257595e+17, 1.278254946357595e+17, 1.278254946457595e+17, 1.278254946557595e+17, 1.278254946657595e+17, 1.278254946757595e+17, 1.278254946857595e+17, 1.278254946957596e+17, 1.278254947057595e+17, 1.278254947157595e+17, 1.278254947257595e+17, 1.278254947357595e+17, 1.278254947457595e+17, 1.278254947557595e+17, 1.278254947657595e+17, 1.278254947757595e+17, 1.278254947857595e+17, 1.278254947957595e+17, 1.278254948057595e+17, 1.278254948157595e+17, 1.278254948257595e+17, 1.278254948357595e+17, 1.278254948457596e+17, 1.278254948557595e+17, 1.278254948657595e+17, 1.278254948757595e+17, 1.278254948857595e+17, 1.278254948957595e+17, 1.278254949057595e+17, 1.278254949157595e+17, 1.278254949257595e+17, 1.278254949357595e+17, 1.278254949457595e+17, 1.278254949557596e+17, 1.278254949657595e+17, 1.278254949757595e+17, 1.278254949857595e+17, 1.278254949957595e+17, 1.278254950057595e+17, 1.278254950157595e+17, 1.278254950257595e+17, 1.278254950357595e+17, 1.278254950457595e+17, 1.278254950557595e+17, 1.278254950657595e+17, 1.278254950757595e+17, 1.278254950857595e+17, 1.278254950957595e+17, 1.278254951057596e+17, 1.278254951157595e+17, 1.278254951257595e+17, 1.278254951357595e+17, 1.278254951457595e+17, 1.278254951557595e+17, 1.278254951657595e+17, 1.278254951757595e+17, 1.278254951857595e+17, 1.278254951957595e+17, 1.278254952057595e+17, 1.278254952157596e+17, 1.278254952257595e+17, 1.278254952357595e+17, 1.278254952457595e+17, 1.278254952557595e+17, 1.278254952657595e+17, 1.278254952757595e+17, 1.278254952857595e+17, 1.278254952957595e+17, 1.278254953057595e+17, 1.278254953157595e+17, 1.278254953257596e+17, 1.278254953357595e+17, 1.278254953457595e+17, 1.278254953557595e+17, 1.278254953657595e+17, 1.278254953757595e+17, 1.278254953857595e+17, 1.278254953957595e+17, 1.278254954057595e+17, 1.278254954157595e+17, 1.278254954257595e+17, 1.278254954357595e+17, 1.278254954457595e+17, 1.278254954557595e+17, 1.278254954657595e+17, 1.278254954757596e+17, 1.278254954857595e+17, 1.278254954957595e+17, 1.278254955057595e+17, 1.278254955157595e+17, 1.278254955257595e+17, 1.278254955357595e+17, 1.278254955457595e+17, 1.278254955557595e+17, 1.278254955657595e+17, 1.278254955757595e+17, 1.278254955857596e+17, 1.278254955957595e+17, 1.278254956057595e+17, 1.278254956157595e+17, 1.278254956257595e+17, 1.278254956357595e+17, 1.278254956457595e+17, 1.278254956557595e+17, 1.278254956657595e+17, 1.278254956757595e+17, 1.278254956857595e+17, 1.278254956957595e+17, 1.278254957057595e+17, 1.278254957157595e+17, 1.278254957257595e+17, 1.278254957357596e+17, 1.278254957457595e+17, 1.278254957557595e+17, 1.278254957657595e+17, 1.278254957757595e+17, 1.278254957857595e+17, 1.278254957957595e+17, 1.278254958057595e+17, 1.278254958157595e+17, 1.278254958257595e+17, 1.278254958357595e+17, 1.278254958457596e+17, 1.278254958557595e+17, 1.278254958657595e+17, 1.278254958757595e+17, 1.278254958857595e+17, 1.278254958957595e+17, 1.278254959057595e+17, 1.278254959157595e+17, 1.278254959257595e+17, 1.278254959357595e+17, 1.278254959457595e+17, 1.278254959557595e+17, 1.278254959657595e+17, 1.278254959757595e+17, 1.278254959857595e+17, 1.278254959957596e+17, 1.278254960057595e+17, 1.278254960157595e+17, 1.278254960257595e+17, 1.278254960357595e+17, 1.278254960457595e+17, 1.278254960557595e+17, 1.278254960657595e+17, 1.278254960757595e+17, 1.278254960857595e+17, 1.278254960957595e+17, 1.278254961057596e+17, 1.278254961157595e+17, 1.278254961257595e+17, 1.278254961357595e+17, 1.278254961457595e+17, 1.278254961557595e+17, 1.278254961657595e+17, 1.278254961757595e+17, 1.278254961857595e+17, 1.278254961957595e+17, 1.278254962057595e+17, 1.278254962157596e+17, 1.278254962257595e+17, 1.278254962357595e+17, 1.278254962457595e+17, 1.278254962557596e+17, 1.278254962657595e+17, 1.278254962757595e+17, 1.278254962857595e+17, 1.278254962957595e+17, 1.278254963057595e+17, 1.278254963157595e+17, 1.278254963257595e+17, 1.278254963357595e+17, 1.278254963457595e+17, 1.278254963557595e+17, 1.278254963657596e+17, 1.278254963757595e+17, 1.278254963857595e+17, 1.278254963957595e+17, 1.278254964057595e+17, 1.278254964157595e+17, 1.278254964257595e+17, 1.278254964357595e+17, 1.278254964457595e+17, 1.278254964557595e+17, 1.278254964657595e+17, 1.278254964757596e+17, 1.278254964857595e+17, 1.278254964957595e+17, 1.278254965057595e+17, 1.278254965157595e+17, 1.278254965257595e+17, 1.278254965357595e+17, 1.278254965457595e+17, 1.278254965557595e+17, 1.278254965657595e+17, 1.278254965757595e+17, 1.278254965857595e+17, 1.278254965957595e+17, 1.278254966057595e+17, 1.278254966157595e+17, 1.278254966257596e+17, 1.278254966357595e+17, 1.278254966457595e+17, 1.278254966557595e+17, 1.278254966657595e+17, 1.278254966757595e+17, 1.278254966857595e+17, 1.278254966957595e+17, 1.278254967057595e+17, 1.278254967157595e+17, 1.278254967257595e+17, 1.278254967357596e+17, 1.278254967457595e+17, 1.278254967557595e+17, 1.278254967657595e+17, 1.278254967757595e+17, 1.278254967857595e+17, 1.278254967957595e+17, 1.278254968057595e+17, 1.278254968157595e+17, 1.278254968257595e+17, 1.278254968357595e+17, 1.278254968457595e+17, 1.278254968557595e+17, 1.278254968657595e+17, 1.278254968757595e+17, 1.278254968857596e+17, 1.278254968957595e+17, 1.278254969057595e+17, 1.278254969157595e+17, 1.278254969257595e+17, 1.278254969357595e+17, 1.278254969457595e+17, 1.278254969557595e+17, 1.278254969657595e+17, 1.278254969757595e+17, 1.278254969857595e+17, 1.278254969957596e+17, 1.278254970057595e+17, 1.278254970157595e+17, 1.278254970257595e+17, 1.278254970357595e+17, 1.278254970457595e+17, 1.278254970557595e+17, 1.278254970657595e+17, 1.278254970757595e+17, 1.278254970857595e+17, 1.278254970957595e+17, 1.278254971057596e+17, 1.278254971157595e+17, 1.278254971257595e+17, 1.278254971357595e+17, 1.278254971457596e+17, 1.278254971557595e+17, 1.278254971657595e+17, 1.278254971757595e+17, 1.278254971857595e+17, 1.278254971957595e+17, 1.278254972057595e+17, 1.278254972157595e+17, 1.278254972257595e+17, 1.278254972357595e+17, 1.278254972457595e+17, 1.278254972557596e+17, 1.278254972657595e+17, 1.278254972757595e+17, 1.278254972857595e+17, 1.278254972957595e+17, 1.278254973057595e+17, 1.278254973157595e+17, 1.278254973257595e+17, 1.278254973357595e+17, 1.278254973457595e+17, 1.278254973557595e+17, 1.278254973657596e+17, 1.278254973757595e+17, 1.278254973857595e+17, 1.278254973957595e+17, 1.278254974057595e+17, 1.278254974157595e+17, 1.278254974257595e+17, 1.278254974357595e+17, 1.278254974457595e+17, 1.278254974557595e+17, 1.278254974657595e+17, 1.278254974757595e+17, 1.278254974857595e+17, 1.278254974957595e+17, 1.278254975057595e+17, 1.278254975157596e+17, 1.278254975257595e+17, 1.278254975357595e+17, 1.278254975457595e+17, 1.278254975557595e+17, 1.278254975657595e+17, 1.278254975757595e+17, 1.278254975857595e+17, 1.278254975957595e+17, 1.278254976057595e+17, 1.278254976157595e+17, 1.278254976257596e+17, 1.278254976357595e+17, 1.278254976457595e+17, 1.278254976557595e+17, 1.278254976657595e+17, 1.278254976757595e+17, 1.278254976857595e+17, 1.278254976957595e+17, 1.278254977057595e+17, 1.278254977157595e+17, 1.278254977257595e+17, 1.278254977357595e+17, 1.278254977457595e+17, 1.278254977557595e+17, 1.278254977657595e+17, 1.278254977757596e+17, 1.278254977857595e+17, 1.278254977957595e+17, 1.278254978057595e+17, 1.278254978157595e+17, 1.278254978257595e+17, 1.278254978357595e+17, 1.278254978457595e+17, 1.278254978557595e+17, 1.278254978657595e+17, 1.278254978757595e+17, 1.278254978857596e+17, 1.278254978957595e+17, 1.278254979057595e+17, 1.278254979157595e+17, 1.278254979257595e+17, 1.278254979357595e+17, 1.278254979457595e+17, 1.278254979557595e+17, 1.278254979657595e+17, 1.278254979757595e+17, 1.278254979857595e+17, 1.278254979957595e+17, 1.278254980057595e+17, 1.278254980157595e+17, 1.278254980257595e+17, 1.278254980357596e+17, 1.278254980457595e+17, 1.278254980557595e+17, 1.278254980657595e+17, 1.278254980757595e+17, 1.278254980857595e+17, 1.278254980957595e+17, 1.278254981057595e+17, 1.278254981157595e+17, 1.278254981257595e+17, 1.278254981357595e+17, 1.278254981457596e+17, 1.278254981557595e+17, 1.278254981657595e+17, 1.278254981757595e+17, 1.278254981857595e+17, 1.278254981957595e+17, 1.278254982057595e+17, 1.278254982157595e+17, 1.278254982257595e+17, 1.278254982357595e+17, 1.278254982457595e+17, 1.278254982557596e+17, 1.278254982657595e+17, 1.278254982757595e+17, 1.278254982857595e+17, 1.278254982957595e+17, 1.278254983057595e+17, 1.278254983157595e+17, 1.278254983257595e+17, 1.278254983357595e+17, 1.278254983457595e+17, 1.278254983557595e+17, 1.278254983657595e+17, 1.278254983757595e+17, 1.278254983857595e+17, 1.278254983957595e+17, 1.278254984057596e+17, 1.278254984157595e+17, 1.278254984257595e+17, 1.278254984357595e+17, 1.278254984457595e+17, 1.278254984557595e+17, 1.278254984657595e+17, 1.278254984757595e+17, 1.278254984857595e+17, 1.278254984957595e+17, 1.278254985057595e+17, 1.278254985157596e+17, 1.278254985257595e+17, 1.278254985357595e+17, 1.278254985457595e+17, 1.278254985557595e+17, 1.278254985657595e+17, 1.278254985757595e+17, 1.278254985857595e+17, 1.278254985957595e+17, 1.278254986057595e+17, 1.278254986157595e+17, 1.278254986257595e+17, 1.278254986357595e+17, 1.278254986457595e+17, 1.278254986557595e+17, 1.278254986657596e+17, 1.278254986757595e+17, 1.278254986857595e+17, 1.278254986957595e+17, 1.278254987057595e+17, 1.278254987157595e+17, 1.278254987257595e+17, 1.278254987357595e+17, 1.278254987457595e+17, 1.278254987557595e+17, 1.278254987657595e+17, 1.278254987757596e+17, 1.278254987857595e+17, 1.278254987957595e+17, 1.278254988057595e+17, 1.278254988157595e+17, 1.278254988257595e+17, 1.278254988357595e+17, 1.278254988457595e+17, 1.278254988557595e+17, 1.278254988657595e+17, 1.278254988757595e+17, 1.278254988857595e+17, 1.278254988957595e+17, 1.278254989057595e+17, 1.278254989157595e+17, 1.278254989257596e+17, 1.278254989357595e+17, 1.278254989457595e+17, 1.278254989557595e+17, 1.278254989657595e+17, 1.278254989757595e+17, 1.278254989857595e+17, 1.278254989957595e+17, 1.278254990057595e+17, 1.278254990157595e+17, 1.278254990257595e+17, 1.278254990357596e+17, 1.278254990457595e+17, 1.278254990557595e+17, 1.278254990657595e+17, 1.278254990757595e+17, 1.278254990857595e+17, 1.278254990957595e+17, 1.278254991057595e+17, 1.278254991157595e+17, 1.278254991257595e+17, 1.278254991357595e+17, 1.278254991457596e+17, 1.278254991557595e+17, 1.278254991657595e+17, 1.278254991757595e+17, 1.278254991857595e+17, 1.278254991957595e+17, 1.278254992057595e+17, 1.278254992157595e+17, 1.278254992257595e+17, 1.278254992357595e+17, 1.278254992457595e+17, 1.278254992557595e+17, 1.278254992657595e+17, 1.278254992757595e+17, 1.278254992857595e+17, 1.278254992957596e+17, 1.278254993057595e+17, 1.278254993157595e+17, 1.278254993257595e+17, 1.278254993357595e+17, 1.278254993457595e+17, 1.278254993557595e+17, 1.278254993657595e+17, 1.278254993757595e+17, 1.278254993857595e+17, 1.278254993957595e+17, 1.278254994057596e+17, 1.278254994157595e+17, 1.278254994257595e+17, 1.278254994357595e+17, 1.278254994457595e+17, 1.278254994557595e+17, 1.278254994657595e+17, 1.278254994757595e+17, 1.278254994857595e+17, 1.278254994957595e+17, 1.278254995057595e+17, 1.278254995157595e+17, 1.278254995257595e+17, 1.278254995357595e+17, 1.278254995457595e+17, 1.278254995557596e+17, 1.278254995657595e+17, 1.278254995757595e+17, 1.278254995857595e+17, 1.278254995957595e+17, 1.278254996057595e+17, 1.278254996157595e+17, 1.278254996257595e+17, 1.278254996357595e+17, 1.278254996457595e+17, 1.278254996557595e+17, 1.278254996657596e+17, 1.278254996757595e+17, 1.278254996857595e+17, 1.278254996957595e+17, 1.278254997057595e+17, 1.278254997157595e+17, 1.278254997257595e+17, 1.278254997357595e+17, 1.278254997457595e+17, 1.278254997557595e+17, 1.278254997657595e+17, 1.278254997757595e+17, 1.278254997857595e+17, 1.278254997957595e+17, 1.278254998057595e+17, 1.278254998157596e+17, 1.278254998257595e+17, 1.278254998357595e+17, 1.278254998457595e+17, 1.278254998557595e+17, 1.278254998657595e+17, 1.278254998757595e+17, 1.278254998857595e+17, 1.278254998957595e+17, 1.278254999057595e+17, 1.278254999157595e+17, 1.278254999257596e+17, 1.278254999357595e+17, 1.278254999457595e+17, 1.278254999557595e+17, 1.278254999657595e+17, 1.278254999757595e+17, 1.278254999857595e+17, 1.278254999957595e+17, 1.278255000057595e+17, 1.278255000157595e+17, 1.278255000257595e+17, 1.278255000357596e+17, 1.278255000457595e+17, 1.278255000557595e+17, 1.278255000657595e+17, 1.278255000757596e+17, 1.278255000857595e+17, 1.278255000957595e+17, 1.278255001057595e+17, 1.278255001157595e+17, 1.278255001257595e+17, 1.278255001357595e+17, 1.278255001457595e+17, 1.278255001557595e+17, 1.278255001657595e+17, 1.278255001757595e+17, 1.278255001857596e+17, 1.278255001957595e+17, 1.278255002057595e+17, 1.278255002157595e+17, 1.278255002257595e+17, 1.278255002357595e+17, 1.278255002457595e+17, 1.278255002557595e+17, 1.278255002657595e+17, 1.278255002757595e+17, 1.278255002857595e+17, 1.278255002957596e+17, 1.278255003057595e+17, 1.278255003157595e+17, 1.278255003257595e+17, 1.278255003357595e+17, 1.278255003457595e+17, 1.278255003557595e+17, 1.278255003657595e+17, 1.278255003757595e+17, 1.278255003857595e+17, 1.278255003957595e+17, 1.278255004057595e+17, 1.278255004157595e+17, 1.278255004257595e+17, 1.278255004357595e+17, 1.278255004457596e+17, 1.278255004557595e+17, 1.278255004657595e+17, 1.278255004757595e+17, 1.278255004857595e+17, 1.278255004957595e+17, 1.278255005057595e+17, 1.278255005157595e+17, 1.278255005257595e+17, 1.278255005357595e+17, 1.278255005457595e+17, 1.278255005557596e+17, 1.278255005657595e+17, 1.278255005757595e+17, 1.278255005857595e+17, 1.278255005957595e+17, 1.278255006057595e+17, 1.278255006157595e+17, 1.278255006257595e+17, 1.278255006357595e+17, 1.278255006457595e+17, 1.278255006557595e+17, 1.278255006657595e+17, 1.278255006757595e+17, 1.278255006857595e+17, 1.278255006957595e+17, 1.278255007057596e+17, 1.278255007157595e+17, 1.278255007257595e+17, 1.278255007357595e+17, 1.278255007457595e+17, 1.278255007557595e+17, 1.278255007657595e+17, 1.278255007757595e+17, 1.278255007857595e+17, 1.278255007957595e+17, 1.278255008057595e+17, 1.278255008157596e+17, 1.278255008257595e+17, 1.278255008357595e+17, 1.278255008457595e+17, 1.278255008557595e+17, 1.278255008657595e+17, 1.278255008757595e+17, 1.278255008857595e+17, 1.278255008957595e+17, 1.278255009057595e+17, 1.278255009157595e+17, 1.278255009257596e+17, 1.278255009357595e+17, 1.278255009457595e+17, 1.278255009557595e+17, 1.278255009657596e+17, 1.278255009757595e+17, 1.278255009857595e+17, 1.278255009957595e+17, 1.278255010057595e+17, 1.278255010157595e+17, 1.278255010257595e+17, 1.278255010357595e+17, 1.278255010457595e+17, 1.278255010557595e+17, 1.278255010657595e+17, 1.278255010757596e+17, 1.278255010857595e+17, 1.278255010957595e+17, 1.278255011057595e+17, 1.278255011157595e+17, 1.278255011257595e+17, 1.278255011357595e+17, 1.278255011457595e+17, 1.278255011557595e+17, 1.278255011657595e+17, 1.278255011757595e+17, 1.278255011857596e+17, 1.278255011957595e+17, 1.278255012057595e+17, 1.278255012157595e+17, 1.278255012257595e+17, 1.278255012357595e+17, 1.278255012457595e+17, 1.278255012557595e+17, 1.278255012657595e+17, 1.278255012757595e+17, 1.278255012857595e+17, 1.278255012957595e+17, 1.278255013057595e+17, 1.278255013157595e+17, 1.278255013257595e+17, 1.278255013357596e+17, 1.278255013457595e+17, 1.278255013557595e+17, 1.278255013657595e+17, 1.278255013757595e+17, 1.278255013857595e+17, 1.278255013957595e+17, 1.278255014057595e+17, 1.278255014157595e+17, 1.278255014257595e+17, 1.278255014357595e+17, 1.278255014457596e+17, 1.278255014557595e+17, 1.278255014657595e+17, 1.278255014757595e+17, 1.278255014857595e+17, 1.278255014957595e+17, 1.278255015057595e+17, 1.278255015157595e+17, 1.278255015257595e+17, 1.278255015357595e+17, 1.278255015457595e+17, 1.278255015557595e+17, 1.278255015657595e+17, 1.278255015757595e+17, 1.278255015857595e+17, 1.278255015957596e+17, 1.278255016057595e+17, 1.278255016157595e+17, 1.278255016257595e+17, 1.278255016357595e+17, 1.278255016457595e+17, 1.278255016557595e+17, 1.278255016657595e+17, 1.278255016757595e+17, 1.278255016857595e+17, 1.278255016957595e+17, 1.278255017057596e+17, 1.278255017157595e+17, 1.278255017257595e+17, 1.278255017357595e+17, 1.278255017457595e+17, 1.278255017557595e+17, 1.278255017657595e+17, 1.278255017757595e+17, 1.278255017857595e+17, 1.278255017957595e+17, 1.278255018057595e+17, 1.278255018157595e+17, 1.278255018257595e+17, 1.278255018357595e+17, 1.278255018457595e+17, 1.278255018557596e+17, 1.278255018657595e+17, 1.278255018757595e+17, 1.278255018857595e+17, 1.278255018957595e+17, 1.278255019057595e+17, 1.278255019157595e+17, 1.278255019257595e+17, 1.278255019357595e+17, 1.278255019457595e+17, 1.278255019557595e+17, 1.278255019657596e+17, 1.278255019757595e+17, 1.278255019857595e+17, 1.278255019957595e+17, 1.278255020057595e+17, 1.278255020157595e+17, 1.278255020257595e+17, 1.278255020357595e+17, 1.278255020457595e+17, 1.278255020557595e+17, 1.278255020657595e+17, 1.278255020757596e+17, 1.278255020857595e+17, 1.278255020957595e+17, 1.278255021057595e+17, 1.278255021157595e+17, 1.278255021257595e+17, 1.278255021357595e+17, 1.278255021457595e+17, 1.278255021557595e+17, 1.278255021657595e+17, 1.278255021757595e+17, 1.278255021857595e+17, 1.278255021957595e+17, 1.278255022057595e+17, 1.278255022157595e+17, 1.278255022257596e+17, 1.278255022357595e+17, 1.278255022457595e+17, 1.278255022557595e+17, 1.278255022657595e+17, 1.278255022757595e+17, 1.278255022857595e+17, 1.278255022957595e+17, 1.278255023057595e+17, 1.278255023157595e+17, 1.278255023257595e+17, 1.278255023357596e+17, 1.278255023457595e+17, 1.278255023557595e+17, 1.278255023657595e+17, 1.278255023757595e+17, 1.278255023857595e+17, 1.278255023957595e+17, 1.278255024057595e+17, 1.278255024157595e+17, 1.278255024257595e+17, 1.278255024357595e+17, 1.278255024457595e+17, 1.278255024557595e+17, 1.278255024657595e+17, 1.278255024757595e+17, 1.278255024857596e+17, 1.278255024957595e+17, 1.278255025057595e+17, 1.278255025157595e+17, 1.278255025257595e+17, 1.278255025357595e+17, 1.278255025457595e+17, 1.278255025557595e+17, 1.278255025657595e+17, 1.278255025757595e+17, 1.278255025857595e+17, 1.278255025957596e+17, 1.278255026057595e+17, 1.278255026157595e+17, 1.278255026257595e+17, 1.278255026357595e+17, 1.278255026457595e+17, 1.278255026557595e+17, 1.278255026657595e+17, 1.278255026757595e+17, 1.278255026857595e+17, 1.278255026957595e+17, 1.278255027057595e+17, 1.278255027157595e+17, 1.278255027257595e+17, 1.278255027357595e+17, 1.278255027457596e+17, 1.278255027557595e+17, 1.278255027657595e+17, 1.278255027757595e+17, 1.278255027857595e+17, 1.278255027957595e+17, 1.278255028057595e+17, 1.278255028157595e+17, 1.278255028257595e+17, 1.278255028357595e+17, 1.278255028457595e+17, 1.278255028557596e+17, 1.278255028657595e+17, 1.278255028757595e+17, 1.278255028857595e+17, 1.278255028957595e+17, 1.278255029057595e+17, 1.278255029157595e+17, 1.278255029257595e+17, 1.278255029357595e+17, 1.278255029457595e+17, 1.278255029557595e+17, 1.278255029657596e+17, 1.278255029757595e+17, 1.278255029857595e+17, 1.278255029957595e+17, 1.278255030057596e+17, 1.278255030157595e+17, 1.278255030257595e+17, 1.278255030357595e+17, 1.278255030457595e+17, 1.278255030557595e+17, 1.278255030657595e+17, 1.278255030757595e+17, 1.278255030857595e+17, 1.278255030957595e+17, 1.278255031057595e+17, 1.278255031157596e+17, 1.278255031257595e+17, 1.278255031357595e+17, 1.278255031457595e+17, 1.278255031557595e+17, 1.278255031657595e+17, 1.278255031757595e+17, 1.278255031857595e+17, 1.278255031957595e+17, 1.278255032057595e+17, 1.278255032157595e+17, 1.278255032257596e+17, 1.278255032357595e+17, 1.278255032457595e+17, 1.278255032557595e+17, 1.278255032657595e+17, 1.278255032757595e+17, 1.278255032857595e+17, 1.278255032957595e+17, 1.278255033057595e+17, 1.278255033157595e+17, 1.278255033257595e+17, 1.278255033357595e+17, 1.278255033457595e+17, 1.278255033557595e+17, 1.278255033657595e+17, 1.278255033757596e+17, 1.278255033857595e+17, 1.278255033957595e+17, 1.278255034057595e+17, 1.278255034157595e+17, 1.278255034257595e+17, 1.278255034357595e+17, 1.278255034457595e+17, 1.278255034557595e+17, 1.278255034657595e+17, 1.278255034757595e+17, 1.278255034857596e+17, 1.278255034957595e+17, 1.278255035057595e+17, 1.278255035157595e+17, 1.278255035257595e+17, 1.278255035357595e+17, 1.278255035457595e+17, 1.278255035557595e+17, 1.278255035657595e+17, 1.278255035757595e+17, 1.278255035857595e+17, 1.278255035957595e+17, 1.278255036057595e+17, 1.278255036157595e+17, 1.278255036257595e+17, 1.278255036357596e+17, 1.278255036457595e+17, 1.278255036557595e+17, 1.278255036657595e+17, 1.278255036757595e+17, 1.278255036857595e+17, 1.278255036957595e+17, 1.278255037057595e+17, 1.278255037157595e+17, 1.278255037257595e+17, 1.278255037357595e+17, 1.278255037457596e+17, 1.278255037557595e+17, 1.278255037657595e+17, 1.278255037757595e+17, 1.278255037857595e+17, 1.278255037957595e+17, 1.278255038057595e+17, 1.278255038157595e+17, 1.278255038257595e+17, 1.278255038357595e+17, 1.278255038457595e+17, 1.278255038557596e+17, 1.278255038657595e+17, 1.278255038757595e+17, 1.278255038857595e+17, 1.278255038957596e+17, 1.278255039057595e+17, 1.278255039157595e+17, 1.278255039257595e+17, 1.278255039357595e+17, 1.278255039457595e+17, 1.278255039557595e+17, 1.278255039657595e+17, 1.278255039757595e+17, 1.278255039857595e+17, 1.278255039957595e+17, 1.278255040057596e+17, 1.278255040157595e+17, 1.278255040257595e+17, 1.278255040357595e+17, 1.278255040457595e+17, 1.278255040557595e+17, 1.278255040657595e+17, 1.278255040757595e+17, 1.278255040857595e+17, 1.278255040957595e+17, 1.278255041057595e+17, 1.278255041157596e+17, 1.278255041257595e+17, 1.278255041357595e+17, 1.278255041457595e+17, 1.278255041557595e+17, 1.278255041657595e+17, 1.278255041757595e+17, 1.278255041857595e+17, 1.278255041957595e+17, 1.278255042057595e+17, 1.278255042157595e+17, 1.278255042257595e+17, 1.278255042357595e+17, 1.278255042457595e+17, 1.278255042557595e+17, 1.278255042657596e+17, 1.278255042757595e+17, 1.278255042857595e+17, 1.278255042957595e+17, 1.278255043057595e+17, 1.278255043157595e+17, 1.278255043257595e+17, 1.278255043357595e+17, 1.278255043457595e+17, 1.278255043557595e+17, 1.278255043657595e+17, 1.278255043757596e+17, 1.278255043857595e+17, 1.278255043957595e+17, 1.278255044057595e+17, 1.278255044157595e+17, 1.278255044257595e+17, 1.278255044357595e+17, 1.278255044457595e+17, 1.278255044557595e+17, 1.278255044657595e+17, 1.278255044757595e+17, 1.278255044857595e+17, 1.278255044957595e+17, 1.278255045057595e+17, 1.278255045157595e+17, 1.278255045257596e+17, 1.278255045357595e+17, 1.278255045457595e+17, 1.278255045557595e+17, 1.278255045657595e+17, 1.278255045757595e+17, 1.278255045857595e+17, 1.278255045957595e+17, 1.278255046057595e+17, 1.278255046157595e+17, 1.278255046257595e+17, 1.278255046357596e+17, 1.278255046457595e+17, 1.278255046557595e+17, 1.278255046657595e+17, 1.278255046757595e+17, 1.278255046857595e+17, 1.278255046957595e+17, 1.278255047057595e+17, 1.278255047157595e+17, 1.278255047257595e+17, 1.278255047357595e+17, 1.278255047457595e+17, 1.278255047557595e+17, 1.278255047657595e+17, 1.278255047757595e+17, 1.278255047857596e+17, 1.278255047957595e+17, 1.278255048057595e+17, 1.278255048157595e+17, 1.278255048257595e+17, 1.278255048357595e+17, 1.278255048457595e+17, 1.278255048557595e+17, 1.278255048657595e+17, 1.278255048757595e+17, 1.278255048857595e+17, 1.278255048957596e+17, 1.278255049057595e+17, 1.278255049157595e+17, 1.278255049257595e+17, 1.278255049357595e+17, 1.278255049457595e+17, 1.278255049557595e+17, 1.278255049657595e+17, 1.278255049757595e+17, 1.278255049857595e+17, 1.278255049957595e+17, 1.278255050057596e+17, 1.278255050157595e+17, 1.278255050257595e+17, 1.278255050357595e+17, 1.278255050457595e+17, 1.278255050557595e+17, 1.278255050657595e+17, 1.278255050757595e+17, 1.278255050857595e+17, 1.278255050957595e+17, 1.278255051057595e+17, 1.278255051157595e+17, 1.278255051257595e+17, 1.278255051357595e+17, 1.278255051457595e+17, 1.278255051557596e+17, 1.278255051657595e+17, 1.278255051757595e+17, 1.278255051857595e+17, 1.278255051957595e+17, 1.278255052057595e+17, 1.278255052157595e+17, 1.278255052257595e+17, 1.278255052357595e+17, 1.278255052457595e+17, 1.278255052557595e+17, 1.278255052657596e+17, 1.278255052757595e+17, 1.278255052857595e+17, 1.278255052957595e+17, 1.278255053057595e+17, 1.278255053157595e+17, 1.278255053257595e+17, 1.278255053357595e+17, 1.278255053457595e+17, 1.278255053557595e+17, 1.278255053657595e+17, 1.278255053757595e+17, 1.278255053857595e+17, 1.278255053957595e+17, 1.278255054057595e+17, 1.278255054157596e+17, 1.278255054257595e+17, 1.278255054357595e+17, 1.278255054457595e+17, 1.278255054557595e+17, 1.278255054657595e+17, 1.278255054757595e+17, 1.278255054857595e+17, 1.278255054957595e+17, 1.278255055057595e+17, 1.278255055157595e+17, 1.278255055257596e+17, 1.278255055357595e+17, 1.278255055457595e+17, 1.278255055557595e+17, 1.278255055657595e+17, 1.278255055757595e+17, 1.278255055857595e+17, 1.278255055957595e+17, 1.278255056057595e+17, 1.278255056157595e+17, 1.278255056257595e+17, 1.278255056357595e+17, 1.278255056457595e+17, 1.278255056557595e+17, 1.278255056657595e+17, 1.278255056757596e+17, 1.278255056857595e+17, 1.278255056957595e+17, 1.278255057057595e+17, 1.278255057157595e+17, 1.278255057257595e+17, 1.278255057357595e+17, 1.278255057457595e+17, 1.278255057557595e+17, 1.278255057657595e+17, 1.278255057757595e+17, 1.278255057857596e+17, 1.278255057957595e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
