netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 29;
			channels = 6;
			categories = 174;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  11.5, 77.9, 79.2, 64.6, 79.0, 73.3, 80.1, 81.1, 46.5, 76.3, 74.8, 73.5, 79.0, 78.8, 79.0, 80.4, 76.5, 74.5, 79.6, 80.0, 79.7, 78.0, 79.9, 80.4, 72.4, 73.9, 78.7, 79.0, 79.5;
			max_depth =  83.2, 80.5, 80.9, 78.7, 81.4, 82.0, 81.5, 82.7, 53.7, 83.1, 77.7, 75.3, 81.1, 81.2, 80.7, 81.5, 78.2, 76.2, 81.0, 81.1, 81.1, 79.5, 81.1, 80.9, 73.6, 76.3, 80.0, 80.9, 80.8;
			start_time = 130432231980169472, 130432232097982080, 130432232251888256, 130432233157357056, 130432233727513216, 130432234533607040, 130432233935638272, 130432235800481920, 130432254258919424, 130432256195481984, 130432268758294528, 130432270831263232, 130432268648919424, 130432268890950784, 130432237320794496, 130432261229232000, 130432261568919552, 130432261938606976, 130432263681575808, 130432264761107072, 130432264938606976, 130432264945794432, 130432265286107008, 130432263955950720, 130432267766575744, 130432267855481984, 130432270270482048, 130432275282356992, 130432275845638272;
			end_time = 130432285856263296, 130432232143294464, 130432232342513152, 130432233220482048, 130432233772825728, 130432234597044480, 130432233971888256, 130432235827669504, 130432254421731968, 130432256313138304, 130432268913450752, 130432270941575680, 130432268802513152, 130432269031263360, 130432237347825792, 130432261258919552, 130432261605950720, 130432262012513152, 130432263822669568, 130432264909075712, 130432265042044416, 130432265034388352, 130432265367200768, 130432264029388160, 130432267907044480, 130432267959075712, 130432270345325824, 130432275380169472, 130432275913607040;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29;
			region_name = "Layer1","Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21","Layer22","Layer23","Layer24","Layer25","Layer26","Layer27","Layer28";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "0", "0", "0", "0", "0", "0", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "6007", "6007", "6007", "6007", "6007", "6007", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "6007", "6007", "6007", "6007", "6007", "6007", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "6007", "6007", "6007", "6007", "6007", "6007", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63;
			mask_times = {1.304322319801695e+17, 1.304322319890758e+17, 1.304322319981382e+17, 1.304322320072008e+17, 1.304322320162632e+17, 1.304322320253257e+17, 1.304322320343882e+17, 1.304322320434508e+17, 1.30432232052357e+17, 1.304322320615757e+17, 1.304322320706382e+17, 1.30432232079857e+17, 1.304322320889196e+17, 1.304322320979821e+17, 1.304322321070445e+17, 1.30432232116107e+17, 1.304322321251695e+17, 1.304322321342321e+17, 1.304322321432945e+17, 1.304322321522007e+17, 1.304322321612632e+17, 1.304322321704819e+17, 1.304322321795444e+17, 1.30432232188607e+17, 1.304322321976695e+17, 1.304322322065757e+17, 1.304322322157946e+17, 1.304322322248571e+17, 1.304322322337632e+17, 1.304322322428257e+17, 1.304322322518883e+17, 1.304322322609508e+17, 1.304322322700133e+17, 1.304322322790757e+17, 1.304322322881382e+17, 1.304322322972008e+17, 1.304322323062633e+17, 1.30432232315482e+17, 1.304322323243882e+17, 1.304322323334508e+17, 1.304322323425132e+17, 1.304322323515757e+17, 1.304322323606382e+17, 1.304322323697007e+17, 1.304322323787633e+17, 1.304322323876695e+17, 1.30432232396732e+17, 1.304322324057946e+17, 1.30432232414857e+17, 1.304322324239195e+17, 1.30432232432982e+17, 1.304322324420444e+17, 1.304322324509508e+17, 1.304322324600133e+17, 1.304322324690758e+17, 1.304322324781384e+17, 1.304322324872008e+17, 1.304322324962633e+17, 1.304322325051695e+17, 1.304322325142321e+17, 1.304322325232945e+17, 1.30432232532357e+17, 1.304322325414195e+17, 1.30432232550482e+17, 1.304322325595446e+17, 1.30432232568607e+17, 1.304322325776695e+17, 1.304322325865757e+17, 1.304322325957944e+17, 1.30432232604857e+17, 1.304322326139195e+17, 1.30432232622982e+17, 1.304322326320445e+17, 1.304322326411071e+17, 1.304322326501696e+17, 1.30432232659232e+17, 1.304322326682945e+17, 1.304322326772008e+17, 1.304322326864195e+17, 1.304322326953257e+17, 1.304322327043882e+17, 1.304322327136069e+17, 1.304322327226694e+17, 1.304322327318883e+17, 1.304322327409508e+17, 1.304322327500133e+17, 1.304322327590757e+17, 1.304322327681382e+17, 1.304322327773569e+17, 1.304322327862633e+17, 1.304322327953257e+17, 1.304322328043882e+17, 1.304322328134508e+17, 1.304322328225133e+17, 1.304322328315757e+17, 1.304322328406382e+17, 1.304322328497007e+17, 1.304322328587633e+17, 1.304322328678258e+17, 1.304322328768883e+17, 1.304322328857946e+17, 1.304322328948571e+17, 1.304322329039195e+17, 1.30432232912982e+17, 1.304322329220444e+17, 1.304322329311069e+17, 1.304322329401695e+17, 1.30432232949232e+17, 1.304322329582945e+17, 1.304322329672008e+17, 1.304322329762633e+17, 1.304322329853257e+17, 1.304322329943882e+17, 1.304322330034508e+17, 1.304322330125132e+17, 1.304322330215757e+17, 1.304322330306382e+17, 1.304322330395444e+17, 1.304322330487633e+17, 1.304322330578258e+17, 1.30432233066732e+17, 1.304322330759508e+17, 1.30432233084857e+17, 1.304322330939195e+17, 1.30432233102982e+17, 1.304322331120445e+17, 1.304322331211071e+17, 1.304322331300133e+17, 1.304322331390758e+17, 1.304322331482945e+17, 1.304322331573571e+17, 1.304322331664196e+17, 1.304322331753257e+17, 1.304322331843882e+17, 1.304322331934508e+17, 1.304322332025133e+17, 1.304322332114195e+17, 1.30432233220482e+17, 1.304322332295444e+17, 1.30432233238607e+17, 1.304322332476695e+17, 1.304322332567319e+17, 1.304322332656383e+17, 1.304322332747008e+17, 1.304322332837633e+17, 1.304322332928257e+17, 1.304322333018883e+17, 1.304322333109508e+17, 1.304322333200132e+17, 1.304322333290757e+17, 1.30432233337982e+17, 1.304322333470445e+17, 1.304322333562633e+17, 1.304322333651695e+17, 1.304322333742321e+17, 1.304322333832946e+17, 1.30432233392357e+17, 1.304322334014195e+17, 1.304322334104819e+17, 1.304322334195444e+17, 1.30432233428607e+17, 1.304322334376695e+17, 1.30432233446732e+17, 1.304322334557944e+17, 1.304322334647008e+17, 1.304322334737632e+17, 1.304322334828257e+17, 1.304322334918883e+17, 1.304322335009507e+17, 1.304322335100132e+17, 1.304322335190757e+17, 1.304322335281382e+17, 1.304322335372008e+17, 1.304322335462633e+17, 1.304322335553258e+17, 1.304322335643884e+17, 1.304322335734508e+17, 1.304322335825133e+17, 1.304322335915757e+17, 1.304322336006382e+17, 1.304322336097007e+17, 1.304322336187633e+17, 1.304322336278257e+17, 1.304322336370445e+17, 1.304322336459507e+17, 1.304322336550132e+17, 1.304322336642321e+17, 1.304322336732945e+17, 1.304322336822008e+17, 1.304322336912632e+17, 1.304322337003258e+17, 1.304322337093883e+17, 1.304322337184507e+17, 1.304322337275132e+17, 1.304322337365757e+17, 1.304322337454821e+17, 1.304322337545445e+17, 1.304322337637632e+17, 1.304322337728257e+17, 1.304322337818883e+17, 1.304322337909508e+17, 1.304322337998569e+17, 1.304322338089194e+17, 1.30432233817982e+17, 1.304322338270445e+17, 1.30432233836107e+17, 1.304322338451695e+17, 1.304322338540758e+17, 1.304322338632946e+17, 1.30432233872357e+17, 1.304322338814195e+17, 1.304322338904819e+17, 1.304322338995444e+17, 1.30432233908607e+17, 1.304322339175133e+17, 1.304322339265757e+17, 1.304322339356383e+17, 1.304322339447008e+17, 1.304322339537633e+17, 1.304322339628257e+17, 1.304322339718883e+17, 1.304322339809507e+17, 1.304322339900132e+17, 1.304322339989196e+17, 1.30432234007982e+17, 1.304322340170445e+17, 1.30432234026107e+17, 1.304322340351695e+17, 1.304322340440756e+17, 1.304322340531382e+17, 1.30432234062357e+17, 1.304322340714195e+17, 1.304322340806382e+17, 1.304322340897007e+17, 1.304322340987633e+17, 1.304322341078257e+17, 1.304322341168882e+17, 1.304322341257944e+17, 1.304322341348571e+17, 1.304322341440758e+17, 1.30432234152982e+17, 1.304322341620445e+17, 1.304322341711069e+17, 1.304322341801695e+17, 1.30432234189232e+17, 1.304322341984507e+17, 1.304322342073571e+17, 1.304322342165757e+17, 1.304322342256383e+17, 1.304322342345445e+17, 1.30432234243607e+17, 1.304322342526696e+17, 1.30432234261732e+17, 1.304322342707945e+17, 1.304322342798569e+17, 1.304322342889194e+17, 1.30432234297982e+17, 1.304322343068883e+17, 1.30432234316107e+17, 1.304322343251695e+17, 1.304322343342321e+17, 1.304322343432945e+17, 1.304322343523571e+17, 1.304322343614195e+17, 1.30432234370482e+17, 1.304322343793883e+17, 1.30432234388607e+17, 1.304322343975132e+17, 1.304322344065757e+17, 1.304322344157944e+17, 1.304322344247008e+17, 1.304322344339195e+17, 1.30432234442982e+17, 1.304322344522007e+17, 1.304322344611071e+17, 1.304322344701696e+17, 1.30432234479232e+17, 1.304322344882945e+17, 1.304322344973569e+17, 1.304322345064195e+17, 1.304322345153257e+17, 1.304322345243882e+17, 1.30432234533607e+17, 1.304322345426694e+17, 1.304322345518883e+17, 1.304322345607945e+17, 1.30432234569857e+17, 1.304322345789196e+17, 1.304322345879821e+17, 1.304322345970445e+17, 1.30432234606107e+17, 1.304322346151695e+17, 1.304322346242319e+17, 1.304322346332945e+17, 1.304322346422008e+17, 1.304322346514195e+17, 1.30432234660482e+17, 1.304322346695444e+17, 1.30432234678607e+17, 1.304322346875132e+17, 1.304322346965756e+17, 1.304322347056383e+17, 1.304322347147007e+17, 1.304322347237632e+17, 1.304322347328257e+17, 1.304322347418883e+17, 1.304322347509508e+17, 1.304322347600133e+17, 1.30432234769232e+17, 1.304322347781382e+17, 1.304322347872008e+17, 1.304322347964196e+17, 1.304322348053257e+17, 1.304322348143882e+17, 1.304322348234508e+17, 1.304322348325133e+17, 1.304322348415757e+17, 1.304322348506382e+17, 1.304322348597007e+17, 1.304322348687633e+17, 1.304322348778258e+17, 1.304322348868883e+17, 1.304322348959507e+17, 1.30432234904857e+17, 1.304322349139195e+17, 1.30432234922982e+17, 1.304322349320445e+17, 1.304322349411071e+17, 1.304322349501696e+17, 1.30432234959232e+17, 1.304322349682945e+17, 1.304322349773571e+17, 1.304322349864195e+17, 1.304322349953257e+17, 1.304322350043882e+17, 1.304322350134508e+17, 1.304322350225133e+17, 1.304322350315758e+17, 1.304322350406383e+17, 1.304322350495444e+17, 1.30432235058607e+17, 1.304322350676695e+17, 1.30432235076732e+17, 1.304322350857944e+17, 1.304322350947008e+17, 1.304322351037633e+17, 1.304322351128257e+17, 1.304322351218883e+17, 1.304322351309507e+17, 1.304322351400132e+17, 1.304322351490757e+17, 1.304322351581382e+17, 1.304322351672008e+17, 1.304322351762633e+17, 1.304322351853258e+17, 1.304322351943884e+17, 1.304322352034508e+17, 1.304322352125133e+17, 1.304322352215758e+17, 1.304322352306382e+17, 1.304322352397007e+17, 1.30432235248607e+17, 1.304322352576695e+17, 1.30432235266732e+17, 1.304322352757946e+17, 1.304322352847007e+17, 1.304322352937632e+17, 1.304322353028257e+17, 1.304322353118883e+17, 1.304322353209508e+17, 1.304322353300132e+17, 1.304322353390757e+17, 1.304322353479821e+17, 1.304322353570445e+17, 1.304322353662633e+17, 1.304322353751694e+17, 1.304322353842319e+17, 1.304322353932945e+17, 1.30432235402357e+17, 1.304322354112632e+17, 1.30432235420482e+17, 1.304322354295446e+17, 1.304322354386071e+17, 1.304322354476695e+17, 1.304322354565757e+17, 1.304322354656383e+17, 1.304322354747008e+17, 1.304322354837632e+17, 1.304322354928257e+17, 1.304322355017321e+17, 1.304322355107945e+17, 1.30432235519857e+17, 1.304322355289194e+17, 1.30432235537982e+17, 1.304322355472008e+17, 1.30432235556107e+17, 1.304322355651695e+17, 1.304322355742319e+17, 1.304322355832945e+17, 1.30432235592357e+17, 1.304322356014195e+17, 1.30432235610482e+17, 1.304322356195446e+17, 1.30432235628607e+17, 1.304322356375132e+17, 1.30432235646732e+17, 1.304322356557944e+17, 1.30432235664857e+17, 1.304322356739195e+17, 1.304322356831382e+17, 1.304322356922007e+17, 1.304322357011071e+17, 1.304322357101695e+17, 1.30432235719232e+17, 1.304322357282945e+17, 1.304322357373571e+17, 1.304322357462632e+17, 1.304322357553257e+17, 1.304322357643882e+17, 1.304322357734508e+17, 1.304322357825133e+17, 1.304322357914195e+17, 1.304322358004819e+17, 1.304322358095444e+17, 1.30432235818607e+17, 1.304322358276695e+17, 1.30432235836732e+17, 1.304322358457944e+17, 1.304322358548571e+17, 1.304322358639195e+17, 1.30432235872982e+17, 1.304322358820445e+17, 1.304322358912632e+17, 1.304322359003258e+17, 1.304322359093883e+17, 1.304322359184508e+17, 1.304322359275132e+17, 1.304322359365757e+17, 1.304322359456383e+17, 1.304322359547007e+17, 1.304322359637632e+17, 1.304322359726696e+17, 1.304322359818883e+17, 1.304322359907945e+17, 1.30432235999857e+17, 1.304322360089196e+17, 1.30432236017982e+17, 1.304322360270445e+17, 1.30432236036107e+17, 1.304322360450132e+17, 1.304322360540758e+17, 1.304322360631383e+17, 1.304322360722008e+17, 1.304322360812632e+17, 1.304322360903258e+17, 1.304322360993883e+17, 1.304322361082944e+17, 1.304322361173569e+17, 1.304322361264195e+17, 1.30432236135482e+17, 1.304322361445445e+17, 1.304322361534508e+17, 1.304322361626696e+17, 1.304322361715757e+17, 1.304322361806382e+17, 1.30432236189857e+17, 1.304322361987633e+17, 1.304322362078258e+17, 1.304322362168883e+17, 1.304322362259508e+17, 1.304322362350132e+17, 1.304322362439195e+17, 1.30432236252982e+17, 1.304322362622007e+17, 1.304322362712632e+17, 1.304322362803256e+17, 1.304322362893882e+17, 1.304322362984507e+17, 1.304322363075132e+17, 1.304322363165757e+17, 1.304322363256383e+17, 1.304322363347008e+17, 1.304322363437633e+17, 1.304322363526694e+17, 1.30432236361732e+17, 1.304322363707945e+17, 1.30432236379857e+17, 1.304322363889196e+17, 1.304322363978258e+17, 1.304322364068883e+17, 1.304322364159507e+17, 1.304322364250132e+17, 1.304322364340756e+17, 1.304322364431382e+17, 1.304322364520445e+17, 1.304322364612632e+17, 1.304322364703258e+17, 1.304322364793883e+17, 1.304322364884508e+17, 1.304322364973571e+17, 1.304322365064195e+17, 1.30432236515482e+17, 1.304322365245444e+17, 1.304322365336069e+17, 1.304322365425133e+17, 1.304322365515757e+17, 1.304322365607945e+17, 1.30432236569857e+17, 1.304322365789196e+17, 1.304322365878258e+17, 1.304322365968882e+17, 1.304322366059507e+17, 1.304322366150132e+17, 1.304322366240758e+17, 1.304322366331383e+17, 1.304322366420445e+17, 1.304322366511071e+17, 1.304322366601695e+17, 1.30432236669232e+17, 1.304322366782944e+17, 1.304322366873569e+17, 1.304322366962633e+17, 1.30432236705482e+17, 1.304322367143884e+17, 1.304322367234508e+17, 1.304322367325133e+17, 1.304322367415758e+17, 1.304322367506382e+17, 1.304322367597007e+17, 1.304322367687633e+17, 1.304322367776695e+17, 1.30432236786732e+17, 1.304322367957944e+17, 1.304322368048571e+17, 1.304322368137632e+17, 1.304322368228257e+17, 1.304322368318883e+17, 1.304322368409508e+17, 1.304322368500132e+17, 1.304322368590757e+17, 1.304322368679821e+17, 1.304322368770445e+17, 1.304322368862633e+17, 1.304322368951694e+17, 1.304322369042319e+17, 1.304322369132945e+17, 1.30432236922357e+17, 1.304322369314195e+17, 1.304322369406382e+17, 1.304322369495446e+17, 1.304322369586071e+17, 1.304322369676695e+17, 1.30432236976732e+17, 1.304322369857946e+17, 1.30432236994857e+17, 1.304322370039195e+17, 1.304322370129819e+17, 1.304322370220444e+17, 1.304322370309508e+17, 1.304322370401695e+17, 1.304322370490757e+17, 1.304322370581382e+17, 1.304322370673571e+17, 1.304322370762633e+17, 1.304322370853257e+17, 1.304322370943882e+17, 1.304322371034508e+17, 1.304322371125133e+17, 1.304322371215757e+17, 1.304322371306383e+17, 1.304322371397007e+17, 1.304322371487633e+17, 1.304322371578258e+17, 1.304322371668883e+17, 1.304322371759508e+17, 1.304322371851695e+17, 1.304322371940756e+17, 1.304322372031382e+17, 1.304322372122007e+17, 1.304322372212632e+17, 1.304322372303258e+17, 1.304322372393883e+17, 1.304322372484508e+17, 1.304322372575133e+17, 1.304322372665757e+17, 1.304322372756383e+17, 1.304322372845445e+17, 1.30432237293607e+17, 1.304322373026694e+17, 1.30432237311732e+17, 1.304322373207945e+17, 1.304322373297009e+17, 1.304322373387633e+17, 1.304322373478258e+17, 1.304322373568882e+17, 1.304322373659507e+17, 1.304322373748571e+17, 1.304322373839195e+17, 1.30432237392982e+17, 1.304322374020445e+17, 1.304322374111071e+17, 1.304322374201696e+17, 1.30432237429232e+17, 1.304322374382944e+17, 1.304322374473569e+17, 1.304322374564195e+17, 1.30432237465482e+17, 1.304322374743882e+17, 1.304322374834508e+17, 1.304322374925133e+17, 1.304322375015758e+17, 1.304322375106382e+17, 1.304322375197007e+17, 1.304322375287633e+17, 1.304322375378257e+17, 1.304322375468882e+17, 1.30432237556107e+17, 1.304322375650132e+17, 1.304322375740758e+17, 1.304322375831383e+17, 1.304322375922008e+17, 1.304322376012632e+17, 1.304322376103258e+17, 1.304322376193883e+17, 1.304322376284507e+17, 1.304322376373569e+17, 1.304322376464195e+17, 1.304322376556383e+17, 1.304322376647008e+17, 1.304322376737633e+17, 1.304322376826696e+17, 1.304322376917321e+17, 1.304322377007945e+17, 1.30432237709857e+17, 1.304322377189194e+17, 1.30432237727982e+17, 1.304322377368883e+17, 1.304322377459508e+17, 1.304322377551695e+17, 1.304322377640758e+17, 1.304322377732945e+17, 1.30432237782357e+17, 1.304322377912632e+17, 1.304322378003256e+17, 1.304322378093882e+17, 1.304322378184507e+17, 1.304322378275132e+17, 1.304322378364196e+17, 1.30432237845482e+17, 1.304322378545445e+17, 1.30432237863607e+17, 1.304322378726694e+17, 1.304322378815757e+17, 1.304322378906382e+17, 1.304322378997007e+17, 1.304322379087633e+17, 1.304322379178258e+17, 1.304322379268883e+17, 1.304322379359508e+17, 1.304322379450132e+17, 1.304322379540758e+17, 1.304322379631382e+17, 1.304322379720445e+17, 1.304322379811071e+17, 1.304322379901696e+17, 1.30432237999232e+17, 1.304322380082945e+17, 1.304322380173571e+17, 1.304322380262633e+17, 1.30432238035482e+17, 1.304322380443882e+17, 1.304322380534508e+17, 1.304322380625133e+17, 1.304322380715757e+17, 1.304322380806383e+17, 1.304322380897007e+17, 1.304322380987633e+17, 1.304322381076695e+17, 1.30432238116732e+17, 1.304322381257944e+17, 1.304322381350132e+17, 1.304322381440758e+17, 1.304322381532945e+17, 1.304322381622008e+17, 1.304322381714195e+17, 1.304322381803258e+17, 1.304322381893883e+17, 1.304322381984508e+17, 1.304322382075133e+17, 1.304322382165757e+17, 1.30432238225482e+17, 1.304322382345445e+17, 1.30432238243607e+17, 1.304322382526694e+17, 1.30432238261732e+17, 1.304322382706382e+17, 1.304322382797007e+17, 1.304322382887631e+17, 1.304322382978257e+17, 1.304322383068882e+17, 1.304322383157944e+17, 1.30432238324857e+17, 1.304322383340758e+17, 1.30432238342982e+17, 1.304322383520445e+17, 1.304322383611069e+17, 1.304322383701695e+17, 1.30432238379232e+17, 1.304322383881382e+17, 1.304322383972008e+17, 1.304322384064196e+17, 1.304322384153258e+17, 1.304322384243884e+17, 1.304322384334508e+17, 1.304322384425133e+17, 1.304322384515757e+17, 1.30432238460482e+17, 1.304322384695444e+17, 1.304322384786071e+17, 1.304322384876695e+17, 1.30432238496732e+17, 1.304322385057946e+17, 1.30432238514857e+17, 1.304322385239195e+17, 1.304322385331383e+17, 1.304322385420444e+17, 1.304322385511069e+17, 1.304322385601695e+17, 1.30432238569232e+17, 1.304322385782945e+17, 1.304322385873571e+17, 1.304322385964196e+17, 1.304322386054821e+17, 1.304322386143882e+17, 1.304322386234508e+17, 1.304322386326694e+17, 1.304322386415757e+17, 1.304322386506382e+17, 1.30432238659857e+17, 1.304322386687633e+17, 1.304322386778258e+17, 1.304322386868883e+17, 1.304322386959508e+17, 1.304322387050132e+17, 1.304322387140758e+17, 1.304322387231382e+17, 1.304322387322007e+17, 1.304322387412632e+17, 1.304322387503258e+17, 1.304322387593883e+17, 1.304322387684508e+17, 1.304322387773571e+17, 1.304322387864195e+17, 1.30432238795482e+17, 1.304322388045445e+17, 1.30432238813607e+17, 1.304322388226694e+17, 1.30432238831732e+17, 1.304322388407945e+17, 1.30432238849857e+17, 1.304322388589196e+17, 1.304322388678258e+17, 1.304322388768882e+17, 1.30432238886107e+17, 1.304322388951695e+17, 1.304322389040756e+17, 1.304322389131382e+17, 1.304322389222007e+17, 1.304322389312632e+17, 1.304322389403258e+17, 1.304322389495444e+17, 1.30432238958607e+17, 1.304322389676695e+17, 1.304322389765757e+17, 1.304322389856383e+17, 1.304322389947007e+17, 1.304322390037632e+17, 1.304322390128257e+17, 1.304322390218883e+17, 1.304322390307945e+17, 1.30432239039857e+17, 1.304322390489196e+17, 1.304322390579821e+17, 1.304322390668882e+17, 1.304322390759507e+17, 1.304322390850132e+17, 1.304322390940758e+17, 1.304322391031383e+17, 1.304322391122008e+17, 1.304322391212632e+17, 1.304322391303258e+17, 1.30432239139232e+17, 1.304322391482944e+17, 1.304322391575132e+17, 1.304322391664195e+17, 1.30432239175482e+17, 1.304322391845445e+17, 1.30432239193607e+17, 1.304322392026696e+17, 1.304322392117321e+17, 1.304322392207945e+17, 1.30432239229857e+17, 1.304322392387633e+17, 1.304322392478258e+17, 1.304322392568883e+17, 1.304322392659508e+17, 1.304322392750132e+17, 1.304322392840758e+17, 1.304322392931383e+17, 1.304322393022008e+17, 1.304322393111069e+17, 1.304322393201695e+17, 1.304322393293882e+17, 1.304322393382945e+17, 1.304322393473571e+17, 1.304322393564195e+17, 1.30432239365482e+17, 1.304322393745445e+17, 1.30432239383607e+17, 1.304322393925133e+17, 1.30432239401732e+17, 1.304322394106382e+17, 1.304322394197007e+17, 1.304322394287633e+17, 1.304322394378258e+17, 1.304322394468883e+17, 1.304322394559508e+17, 1.304322394650132e+17, 1.304322394739195e+17, 1.30432239482982e+17, 1.304322394920445e+17, 1.304322395011071e+17, 1.304322395101696e+17, 1.30432239519232e+17, 1.304322395282945e+17, 1.304322395373571e+17, 1.304322395462633e+17, 1.304322395553257e+17, 1.304322395643882e+17, 1.304322395734508e+17, 1.304322395825133e+17, 1.304322395915757e+17, 1.304322396006382e+17, 1.304322396097007e+17, 1.304322396187633e+17, 1.304322396278258e+17, 1.304322396367319e+17, 1.304322396457944e+17, 1.30432239654857e+17, 1.304322396639195e+17, 1.30432239672982e+17, 1.304322396818883e+17, 1.304322396909508e+17, 1.304322397000132e+17, 1.304322397090757e+17, 1.304322397181382e+17, 1.304322397270445e+17, 1.30432239736107e+17, 1.304322397451695e+17, 1.304322397542321e+17, 1.304322397632945e+17, 1.30432239772357e+17, 1.304322397812632e+17, 1.30432239790482e+17, 1.304322397995444e+17, 1.30432239808607e+17, 1.304322398176695e+17, 1.30432239826732e+17, 1.304322398356383e+17, 1.304322398447008e+17, 1.304322398537632e+17, 1.304322398628257e+17, 1.304322398718883e+17, 1.304322398809507e+17, 1.304322398900132e+17, 1.304322398990757e+17, 1.304322399081382e+17, 1.304322399172008e+17, 1.30432239926107e+17, 1.304322399351695e+17, 1.304322399442319e+17, 1.304322399532945e+17, 1.30432239962357e+17, 1.304322399714195e+17, 1.304322399803258e+17, 1.304322399895444e+17, 1.30432239998607e+17, 1.304322400076695e+17, 1.304322400165757e+17, 1.304322400256383e+17, 1.304322400347008e+17, 1.304322400437632e+17, 1.304322400528257e+17, 1.304322400618883e+17, 1.304322400709508e+17, 1.304322400800133e+17, 1.304322400890757e+17, 1.30432240097982e+17, 1.304322401070445e+17, 1.30432240116107e+17, 1.304322401251694e+17, 1.304322401342319e+17, 1.304322401432945e+17, 1.304322401522008e+17, 1.304322401614195e+17, 1.30432240170482e+17, 1.304322401793883e+17, 1.304322401886071e+17, 1.304322401976695e+17, 1.30432240206732e+17, 1.304322402156383e+17, 1.304322402247008e+17, 1.304322402337633e+17, 1.304322402428257e+17, 1.304322402518883e+17, 1.304322402609508e+17, 1.304322402700133e+17, 1.304322402789194e+17, 1.304322402882945e+17, 1.304322402973571e+17, 1.304322403064196e+17, 1.304322403153257e+17, 1.304322403243882e+17, 1.304322403334508e+17, 1.304322403425133e+17, 1.304322403515758e+17, 1.304322403606383e+17, 1.304322403697009e+17, 1.304322403787633e+17, 1.304322403878258e+17, 1.304322403968882e+17, 1.304322404059507e+17, 1.30432240414857e+17, 1.304322404239195e+17, 1.30432240432982e+17, 1.304322404420445e+17, 1.304322404511071e+17, 1.304322404601696e+17, 1.30432240469232e+17, 1.304322404781382e+17, 1.304322404872008e+17, 1.304322404962633e+17, 1.30432240505482e+17, 1.304322405143882e+17, 1.304322405234508e+17, 1.304322405325133e+17, 1.304322405415758e+17, 1.304322405506383e+17, 1.304322405597007e+17, 1.304322405687633e+17, 1.304322405776695e+17, 1.30432240586732e+17, 1.304322405957946e+17, 1.304322406048571e+17, 1.304322406137632e+17, 1.304322406228257e+17, 1.304322406318883e+17, 1.304322406409508e+17, 1.304322406500133e+17, 1.304322406590757e+17, 1.304322406679821e+17, 1.304322406770446e+17, 1.30432240686107e+17, 1.304322406951695e+17, 1.304322407042319e+17, 1.304322407132945e+17, 1.30432240722357e+17, 1.304322407314195e+17, 1.304322407403258e+17, 1.304322407493883e+17, 1.30432240758607e+17, 1.304322407676695e+17, 1.304322407765757e+17, 1.304322407857946e+17, 1.304322407948571e+17, 1.304322408039195e+17, 1.304322408128257e+17, 1.304322408218883e+17, 1.304322408309508e+17, 1.304322408400133e+17, 1.304322408490757e+17, 1.304322408581384e+17, 1.304322408672008e+17, 1.304322408762633e+17, 1.304322408853257e+17, 1.304322408942321e+17, 1.304322409034508e+17, 1.304322409125132e+17, 1.304322409214195e+17, 1.30432240930482e+17, 1.304322409395444e+17, 1.30432240948607e+17, 1.304322409576695e+17, 1.30432240966732e+17, 1.304322409757944e+17, 1.30432240984857e+17, 1.304322409939195e+17, 1.304322410031382e+17, 1.304322410122007e+17, 1.304322410212632e+17, 1.304322410301695e+17, 1.30432241039232e+17, 1.304322410482945e+17, 1.304322410573571e+17, 1.304322410664196e+17, 1.30432241075482e+17, 1.304322410845445e+17, 1.304322410936069e+17, 1.304322411026694e+17, 1.304322411115757e+17, 1.304322411207945e+17, 1.30432241129857e+17, 1.304322411387633e+17, 1.304322411478258e+17, 1.304322411568882e+17, 1.304322411659507e+17, 1.304322411750132e+17, 1.304322411840758e+17, 1.304322411931383e+17, 1.304322412022007e+17, 1.304322412112632e+17, 1.304322412203258e+17, 1.304322412293883e+17, 1.304322412382945e+17, 1.304322412473569e+17, 1.304322412564195e+17, 1.30432241265482e+17, 1.304322412745444e+17, 1.30432241283607e+17, 1.304322412926694e+17, 1.30432241301732e+17, 1.304322413107945e+17, 1.30432241319857e+17, 1.304322413287633e+17, 1.304322413378257e+17, 1.304322413468882e+17, 1.304322413559507e+17, 1.304322413650132e+17, 1.304322413740758e+17, 1.304322413831383e+17, 1.304322413922008e+17, 1.304322414012634e+17, 1.304322414103258e+17, 1.304322414193883e+17, 1.304322414284508e+17, 1.304322414373571e+17, 1.304322414464195e+17, 1.30432241455482e+17, 1.304322414645445e+17, 1.30432241473607e+17, 1.304322414826696e+17, 1.304322414917321e+17, 1.304322415007945e+17, 1.30432241509857e+17, 1.304322415190758e+17, 1.30432241527982e+17, 1.304322415372008e+17, 1.304322415462632e+17, 1.304322415551695e+17, 1.304322415642321e+17, 1.304322415732945e+17, 1.30432241582357e+17, 1.304322415914195e+17, 1.30432241600482e+17, 1.304322416093883e+17, 1.30432241618607e+17, 1.304322416276695e+17, 1.304322416367319e+17, 1.304322416456383e+17, 1.304322416547008e+17, 1.304322416637632e+17, 1.304322416728257e+17, 1.304322416818883e+17, 1.304322416909508e+17, 1.304322417000133e+17, 1.304322417090757e+17, 1.304322417181382e+17, 1.304322417270445e+17, 1.30432241736107e+17, 1.304322417451695e+17, 1.304322417542321e+17, 1.304322417632946e+17, 1.30432241772357e+17, 1.304322417812632e+17, 1.304322417904819e+17, 1.304322417993883e+17, 1.304322418084508e+17, 1.304322418176695e+17, 1.304322418265757e+17, 1.304322418356383e+17, 1.30432241844857e+17, 1.304322418537633e+17, 1.304322418628257e+17, 1.304322418718883e+17, 1.304322418809507e+17, 1.304322418900132e+17, 1.304322418990757e+17, 1.30432241907982e+17, 1.304322419172008e+17, 1.304322419262633e+17, 1.304322419351695e+17, 1.304322419443884e+17, 1.304322419532945e+17, 1.30432241962357e+17, 1.304322419714195e+17, 1.30432241980482e+17, 1.304322419895444e+17, 1.304322419984508e+17, 1.304322420075133e+17, 1.30432242016732e+17, 1.304322420257946e+17, 1.304322420347007e+17, 1.304322420439195e+17, 1.304322420528257e+17, 1.304322420618883e+17, 1.304322420709508e+17, 1.304322420800132e+17, 1.304322420890757e+17, 1.304322420981382e+17, 1.304322421070445e+17, 1.304322421162633e+17, 1.304322421251694e+17, 1.304322421343882e+17, 1.304322421432945e+17, 1.30432242152357e+17, 1.304322421614195e+17, 1.30432242170482e+17, 1.304322421795446e+17, 1.304322421886071e+17, 1.304322421976695e+17, 1.304322422065757e+17, 1.304322422157946e+17, 1.30432242224857e+17, 1.304322422339195e+17, 1.304322422428257e+17, 1.304322422518883e+17, 1.304322422609508e+17, 1.304322422700133e+17, 1.304322422790757e+17, 1.30432242287982e+17, 1.304322422970445e+17, 1.30432242306107e+17, 1.304322423153257e+17, 1.304322423242319e+17, 1.304322423332945e+17, 1.304322423425133e+17, 1.304322423514195e+17, 1.30432242360482e+17, 1.304322423695446e+17, 1.30432242378607e+17, 1.304322423876695e+17, 1.30432242396732e+17, 1.304322424057944e+17, 1.30432242414857e+17, 1.304322424237633e+17, 1.304322424328257e+17, 1.304322424418883e+17, 1.304322424509508e+17, 1.304322424600133e+17, 1.304322424690757e+17, 1.304322424781382e+17, 1.304322424870445e+17, 1.30432242496107e+17, 1.304322425051695e+17, 1.304322425143882e+17, 1.304322425232945e+17, 1.30432242532357e+17, 1.304322425414195e+17, 1.304322425504819e+17, 1.304322425595444e+17, 1.30432242568607e+17, 1.304322425776695e+17, 1.30432242586732e+17, 1.304322425957944e+17, 1.304322426048571e+17, 1.304322426139195e+17, 1.304322426228257e+17, 1.304322426318883e+17, 1.304322426409508e+17, 1.304322426500132e+17, 1.304322426590757e+17, 1.304322426681382e+17, 1.304322426772008e+17, 1.304322426862633e+17, 1.304322426951695e+17, 1.304322427042321e+17, 1.304322427134508e+17, 1.304322427225133e+17, 1.304322427315758e+17, 1.304322427406382e+17, 1.304322427497007e+17, 1.304322427589196e+17, 1.304322427678257e+17, 1.304322427768883e+17, 1.304322427859507e+17, 1.304322427950132e+17, 1.304322428040758e+17, 1.30432242812982e+17, 1.304322428220445e+17, 1.304322428311069e+17, 1.304322428401695e+17, 1.30432242849232e+17, 1.304322428581382e+17, 1.304322428672008e+17, 1.304322428762633e+17, 1.304322428853258e+17, 1.304322428943882e+17, 1.304322429034508e+17, 1.304322429125132e+17, 1.304322429215757e+17, 1.304322429306382e+17, 1.304322429397007e+17, 1.304322429487633e+17, 1.304322429576695e+17, 1.30432242966732e+17, 1.304322429757946e+17, 1.30432242984857e+17, 1.304322429939195e+17, 1.30432243002982e+17, 1.304322430118883e+17, 1.304322430209508e+17, 1.304322430300133e+17, 1.304322430390758e+17, 1.304322430481384e+17, 1.304322430572008e+17, 1.304322430662633e+17, 1.304322430751695e+17, 1.304322430842321e+17, 1.304322430932945e+17, 1.30432243102357e+17, 1.304322431114195e+17, 1.30432243120482e+17, 1.304322431293883e+17, 1.304322431384507e+17, 1.304322431475132e+17, 1.304322431565757e+17, 1.304322431656383e+17, 1.304322431747008e+17, 1.304322431837632e+17, 1.30432243192982e+17, 1.304322432020445e+17, 1.304322432111071e+17, 1.304322432201696e+17, 1.30432243229232e+17, 1.304322432382945e+17, 1.304322432472008e+17, 1.304322432562633e+17, 1.304322432653257e+17, 1.304322432743882e+17, 1.304322432834508e+17, 1.304322432925133e+17, 1.304322433015757e+17, 1.304322433106383e+17, 1.304322433195444e+17, 1.30432243328607e+17, 1.304322433376695e+17, 1.30432243346732e+17, 1.304322433557944e+17, 1.30432243364857e+17, 1.304322433739195e+17, 1.30432243382982e+17, 1.304322433918883e+17, 1.304322434009507e+17, 1.304322434101695e+17, 1.304322434190757e+17, 1.304322434281382e+17, 1.304322434372008e+17, 1.304322434462633e+17, 1.304322434553258e+17, 1.304322434643884e+17, 1.304322434734508e+17, 1.304322434825133e+17, 1.304322434915758e+17, 1.304322435006382e+17, 1.304322435097007e+17, 1.304322435187633e+17, 1.304322435278257e+17, 1.304322435368882e+17, 1.304322435459507e+17, 1.304322435550132e+17, 1.304322435640758e+17, 1.304322435731383e+17, 1.304322435822008e+17, 1.304322435912634e+17, 1.304322436003258e+17, 1.30432243609232e+17, 1.304322436182945e+17, 1.304322436275132e+17, 1.304322436365757e+17, 1.30432243645482e+17, 1.304322436545445e+17, 1.30432243663607e+17, 1.304322436726696e+17, 1.304322436817321e+17, 1.304322436907945e+17, 1.304322436997007e+17, 1.304322437087633e+17, 1.304322437178257e+17, 1.304322437268882e+17, 1.304322437359507e+17, 1.304322437450132e+17, 1.304322437539195e+17, 1.304322437629819e+17, 1.304322437720444e+17, 1.304322437811069e+17, 1.304322437901695e+17, 1.30432243799232e+17, 1.304322438082945e+17, 1.304322438173571e+17, 1.304322438264196e+17, 1.304322438354821e+17, 1.304322438445445e+17, 1.30432243853607e+17, 1.304322438626694e+17, 1.30432243871732e+17, 1.304322438807945e+17, 1.30432243889857e+17, 1.304322438989194e+17, 1.304322439078258e+17, 1.304322439168883e+17, 1.30432243926107e+17, 1.304322439351695e+17, 1.304322439440756e+17, 1.304322439531382e+17, 1.304322439622007e+17, 1.304322439712632e+17, 1.304322439803258e+17, 1.304322439893883e+17, 1.304322439982945e+17, 1.304322440073571e+17, 1.304322440164195e+17, 1.30432244025482e+17, 1.304322440345445e+17, 1.30432244043607e+17, 1.304322440526694e+17, 1.304322440615758e+17, 1.304322440707945e+17, 1.30432244079857e+17, 1.304322440887633e+17, 1.304322440979821e+17, 1.304322441068882e+17, 1.304322441159507e+17, 1.304322441251695e+17, 1.304322441340756e+17, 1.304322441431382e+17, 1.30432244152357e+17, 1.304322441612632e+17, 1.304322441703258e+17, 1.304322441793883e+17, 1.304322441884508e+17, 1.304322441975133e+17, 1.304322442065757e+17, 1.304322442156383e+17, 1.304322442247007e+17, 1.304322442337632e+17, 1.30432244242982e+17, 1.304322442520444e+17, 1.304322442609508e+17, 1.304322442700133e+17, 1.304322442790757e+17, 1.304322442881382e+17, 1.304322442972008e+17, 1.30432244306107e+17, 1.304322443151694e+17, 1.304322443242319e+17, 1.304322443332945e+17, 1.30432244342357e+17, 1.304322443514195e+17, 1.30432244360482e+17, 1.304322443693883e+17, 1.304322443784507e+17, 1.304322443875132e+17, 1.304322443965757e+17, 1.304322444056383e+17, 1.304322444147008e+17, 1.304322444237633e+17, 1.304322444328257e+17, 1.304322444418883e+17, 1.304322444509508e+17, 1.30432244459857e+17, 1.304322444689194e+17, 1.30432244477982e+17, 1.304322444870445e+17, 1.30432244496107e+17, 1.304322445050132e+17, 1.304322445140758e+17, 1.304322445232945e+17, 1.30432244532357e+17, 1.304322445414195e+17, 1.304322445503256e+17, 1.304322445593882e+17, 1.304322445684507e+17, 1.304322445775132e+17, 1.304322445865757e+17, 1.304322445956383e+17, 1.304322446047008e+17, 1.304322446137633e+17, 1.304322446228257e+17, 1.304322446318883e+17, 1.304322446409508e+17, 1.304322446500132e+17, 1.304322446589196e+17, 1.304322446679821e+17, 1.304322446770445e+17, 1.30432244686107e+17, 1.304322446953257e+17, 1.304322447042321e+17, 1.304322447132945e+17, 1.30432244722357e+17, 1.304322447314195e+17, 1.304322447404819e+17, 1.304322447493883e+17, 1.304322447584507e+17, 1.304322447675132e+17, 1.304322447765757e+17, 1.304322447856383e+17, 1.304322447947008e+17, 1.304322448036069e+17, 1.304322448126694e+17, 1.304322448218883e+17, 1.304322448309508e+17, 1.304322448400133e+17, 1.304322448489196e+17, 1.304322448579821e+17, 1.304322448670445e+17, 1.30432244876107e+17, 1.304322448851695e+17, 1.304322448942319e+17, 1.304322449032945e+17, 1.30432244912357e+17, 1.304322449214195e+17, 1.304322449304819e+17, 1.304322449393883e+17, 1.30432244948607e+17, 1.304322449575133e+17, 1.304322449665757e+17, 1.304322449756383e+17, 1.304322449847007e+17, 1.304322449937632e+17, 1.304322450028257e+17, 1.304322450118883e+17, 1.304322450209508e+17, 1.304322450300133e+17, 1.30432245039232e+17, 1.304322450481382e+17, 1.304322450572008e+17, 1.304322450662633e+17, 1.304322450753258e+17, 1.304322450843882e+17, 1.304322450934508e+17, 1.30432245102357e+17, 1.304322451114195e+17, 1.30432245120482e+17, 1.304322451295444e+17, 1.30432245138607e+17, 1.304322451476695e+17, 1.304322451565757e+17, 1.304322451656383e+17, 1.304322451747007e+17, 1.304322451837632e+17, 1.304322451928257e+17, 1.304322452018883e+17, 1.304322452109508e+17, 1.304322452200133e+17, 1.304322452290758e+17, 1.304322452381382e+17, 1.304322452472008e+17, 1.30432245256107e+17, 1.304322452651695e+17, 1.304322452742321e+17, 1.304322452832945e+17, 1.30432245292357e+17, 1.304322453014195e+17, 1.30432245310482e+17, 1.304322453195446e+17, 1.30432245328607e+17, 1.304322453376695e+17, 1.304322453465757e+17, 1.304322453556383e+17, 1.304322453647008e+17, 1.304322453737633e+17, 1.304322453828257e+17, 1.304322453918883e+17, 1.304322454009508e+17, 1.30432245409857e+17, 1.304322454190757e+17, 1.304322454281382e+17, 1.304322454372008e+17, 1.304322454462633e+17, 1.304322454551695e+17, 1.304322454642321e+17, 1.304322454732946e+17, 1.30432245482357e+17, 1.304322454914195e+17, 1.304322455003258e+17, 1.304322455093883e+17, 1.304322455184508e+17, 1.304322455275133e+17, 1.304322455365757e+17, 1.304322455456383e+17, 1.304322455547008e+17, 1.304322455637633e+17, 1.304322455728257e+17, 1.304322455818883e+17, 1.304322455907945e+17, 1.30432245599857e+17, 1.304322456089196e+17, 1.304322456181382e+17, 1.304322456270445e+17, 1.304322456362633e+17, 1.304322456453258e+17, 1.304322456543884e+17, 1.304322456634508e+17, 1.30432245672357e+17, 1.304322456815757e+17, 1.30432245690482e+17, 1.304322456995444e+17, 1.30432245708607e+17, 1.304322457176695e+17, 1.30432245726732e+17, 1.304322457359507e+17, 1.304322457448571e+17, 1.304322457539195e+17, 1.30432245762982e+17, 1.304322457720444e+17, 1.304322457811069e+17, 1.304322457901695e+17, 1.304322457990757e+17, 1.304322458081382e+17, 1.304322458172008e+17, 1.304322458262633e+17, 1.304322458353258e+17, 1.304322458443882e+17, 1.304322458532945e+17, 1.30432245862357e+17, 1.304322458714195e+17, 1.30432245880482e+17, 1.304322458895446e+17, 1.304322458984507e+17, 1.304322459075132e+17, 1.30432245916732e+17, 1.304322459257944e+17, 1.304322459347008e+17, 1.304322459439195e+17, 1.304322459528257e+17, 1.304322459618883e+17, 1.304322459709508e+17, 1.304322459800133e+17, 1.304322459890757e+17, 1.30432245997982e+17, 1.304322460070445e+17, 1.304322460162632e+17, 1.304322460253257e+17, 1.304322460343882e+17, 1.304322460434508e+17, 1.304322460525133e+17, 1.304322460614195e+17, 1.30432246070482e+17, 1.304322460795446e+17, 1.30432246088607e+17, 1.304322460976695e+17, 1.30432246106732e+17, 1.304322461157944e+17, 1.30432246124857e+17, 1.304322461339195e+17, 1.304322461428257e+17, 1.304322461518883e+17, 1.304322461609508e+17, 1.304322461700132e+17, 1.304322461790757e+17, 1.304322461879821e+17, 1.304322461970445e+17, 1.30432246206107e+17, 1.304322462151695e+17, 1.304322462242321e+17, 1.304322462331382e+17, 1.304322462422007e+17, 1.304322462512632e+17, 1.304322462603258e+17, 1.304322462693883e+17, 1.304322462784507e+17, 1.304322462875132e+17, 1.304322462965757e+17, 1.304322463056383e+17, 1.304322463147008e+17, 1.304322463237633e+17, 1.304322463776695e+17, 1.304322463867319e+17, 1.304322463959507e+17, 1.304322464050132e+17, 1.304322464140758e+17, 1.30432246422982e+17, 1.304322464320445e+17, 1.304322464411071e+17, 1.304322464501696e+17, 1.30432246459232e+17, 1.304322464682945e+17, 1.304322464773569e+17, 1.304322464864195e+17, 1.30432246495482e+17, 1.304322465045445e+17, 1.304322465134508e+17, 1.304322465225133e+17, 1.304322465315758e+17, 1.304322465406382e+17, 1.304322465497007e+17, 1.304322465587631e+17, 1.304322465678257e+17, 1.304322465768882e+17, 1.304322465859507e+17, 1.304322465950132e+17, 1.304322466040758e+17, 1.30432246612982e+17, 1.304322466220445e+17, 1.304322466311069e+17, 1.304322466401695e+17, 1.30432246649232e+17, 1.304322466582945e+17, 1.304322466673571e+17, 1.304322466764195e+17, 1.304322466853258e+17, 1.304322466945445e+17, 1.304322467034508e+17, 1.304322467125133e+17, 1.304322467215757e+17, 1.304322467306382e+17, 1.304322467397007e+17, 1.30432246748607e+17, 1.304322467576695e+17, 1.30432246766732e+17, 1.304322467757946e+17, 1.30432246784857e+17, 1.304322467939195e+17, 1.304322468028257e+17, 1.304322468118883e+17, 1.304322468209508e+17, 1.304322468300133e+17, 1.304322468390757e+17, 1.304322468481382e+17, 1.304322468572008e+17, 1.30432246866107e+17, 1.304322468753257e+17, 1.304322468843882e+17, 1.304322468932945e+17, 1.30432246902357e+17, 1.304322469114195e+17, 1.30432246920482e+17, 1.304322469295446e+17, 1.304322469386071e+17, 1.304322469475132e+17, 1.30432246956732e+17, 1.304322469657944e+17, 1.30432246974857e+17, 1.304322469837633e+17, 1.304322469928257e+17, 1.304322470018883e+17, 1.304322470109508e+17, 1.304322470200133e+17, 1.304322470290757e+17, 1.304322470381382e+17, 1.304322470470445e+17, 1.304322470562632e+17, 1.304322470653257e+17, 1.304322470742321e+17, 1.304322470834508e+17, 1.30432247092357e+17, 1.304322471014195e+17, 1.30432247110482e+17, 1.304322471195444e+17, 1.30432247128607e+17, 1.304322471376695e+17, 1.30432247146732e+17, 1.304322471557944e+17, 1.30432247164857e+17, 1.304322471740756e+17, 1.30432247182982e+17, 1.304322471922007e+17, 1.304322472012632e+17, 1.304322472101696e+17, 1.30432247219232e+17, 1.304322472282945e+17, 1.304322472373569e+17, 1.304322472464195e+17, 1.30432247255482e+17, 1.304322472645445e+17, 1.30432247273607e+17, 1.304322472826696e+17, 1.304322472917321e+17, 1.304322473007945e+17, 1.304322473100132e+17, 1.304322473190757e+17, 1.304322473281382e+17, 1.304322473372008e+17, 1.304322473462633e+17, 1.304322473553258e+17, 1.304322473643882e+17, 1.304322473734508e+17, 1.304322473825133e+17, 1.304322473914195e+17, 1.30432247400482e+17, 1.304322474095446e+17, 1.304322474186071e+17, 1.304322474275132e+17, 1.304322474365757e+17, 1.304322474456383e+17, 1.304322474547008e+17, 1.304322474637632e+17, 1.304322474728257e+17, 1.304322474818883e+17, 1.304322474909508e+17, 1.304322475000133e+17, 1.30432247509232e+17, 1.304322475181382e+17, 1.304322475272008e+17, 1.304322475362632e+17, 1.304322475453257e+17, 1.304322475543882e+17, 1.304322475634508e+17, 1.304322475725133e+17, 1.304322475815758e+17, 1.30432247590482e+17, 1.304322475995446e+17, 1.30432247608607e+17, 1.304322476176695e+17, 1.30432247626732e+17, 1.304322476356383e+17, 1.304322476447008e+17, 1.304322476537633e+17, 1.304322476628257e+17, 1.304322476718883e+17, 1.304322476809508e+17, 1.304322476900133e+17, 1.304322476990757e+17, 1.304322477082945e+17, 1.304322477172008e+17, 1.304322477262632e+17, 1.304322477353257e+17, 1.304322477443882e+17, 1.304322477534508e+17, 1.304322477625133e+17, 1.304322477714195e+17, 1.304322477806383e+17, 1.304322477895444e+17, 1.30432247798607e+17, 1.304322478078257e+17, 1.304322478168882e+17, 1.304322478259507e+17, 1.304322478350132e+17, 1.304322478440756e+17, 1.304322478531382e+17, 1.304322478622007e+17, 1.304322478712632e+17, 1.304322478803258e+17, 1.30432247889232e+17, 1.304322478982944e+17, 1.304322479073569e+17, 1.304322479164195e+17, 1.30432247925482e+17, 1.304322479345445e+17, 1.304322479434508e+17, 1.304322479525133e+17, 1.304322479615758e+17, 1.304322479706382e+17, 1.304322479797007e+17, 1.30432247988607e+17, 1.304322479976695e+17, 1.304322480068883e+17, 1.304322480157946e+17, 1.304322480248571e+17, 1.304322480339195e+17, 1.30432248042982e+17, 1.304322480520444e+17, 1.304322480611069e+17, 1.304322480701695e+17, 1.30432248079232e+17, 1.304322480881382e+17, 1.304322480972008e+17, 1.304322481064195e+17, 1.30432248115482e+17, 1.304322481245445e+17, 1.304322481334508e+17, 1.304322481425132e+17, 1.304322481515757e+17, 1.304322481606382e+17, 1.304322481697007e+17, 1.304322481787633e+17, 1.304322481876695e+17, 1.30432248196732e+17, 1.304322482057946e+17, 1.30432248214857e+17, 1.304322482239195e+17, 1.30432248232982e+17, 1.304322482418883e+17, 1.304322482511071e+17, 1.304322482601695e+17, 1.304322482690758e+17, 1.304322482782945e+17, 1.304322482872008e+17, 1.304322482962632e+17, 1.30432248305482e+17, 1.304322483143882e+17, 1.304322483236069e+17, 1.304322483326694e+17, 1.304322483415757e+17, 1.304322483506382e+17, 1.304322483597007e+17, 1.304322483687633e+17, 1.304322483778258e+17, 1.304322483868883e+17, 1.304322483959507e+17, 1.304322484050132e+17, 1.304322484139195e+17, 1.30432248422982e+17, 1.304322484320445e+17, 1.304322484411071e+17, 1.304322484501696e+17, 1.30432248459232e+17, 1.304322484681382e+17, 1.304322484773571e+17, 1.304322484862633e+17, 1.304322484953257e+17, 1.304322485043882e+17, 1.304322485134508e+17, 1.304322485225133e+17, 1.304322485314195e+17, 1.304322485404819e+17, 1.304322485495444e+17, 1.30432248558607e+17, 1.304322485676695e+17, 1.304322485765757e+17, 1.304322485857944e+17, 1.30432248594857e+17, 1.304322486039195e+17, 1.30432248612982e+17, 1.304322486218883e+17, 1.304322486309507e+17, 1.304322486400132e+17, 1.304322486490757e+17, 1.304322486581382e+17, 1.304322486672008e+17, 1.304322486762633e+17, 1.304322486853258e+17, 1.304322486942321e+17, 1.304322487032945e+17, 1.304322487125133e+17, 1.304322487214195e+17, 1.30432248730482e+17, 1.304322487395444e+17, 1.30432248748607e+17, 1.304322487576695e+17, 1.304322487665757e+17, 1.304322487756383e+17, 1.304322487847007e+17, 1.304322487937632e+17, 1.304322488028257e+17, 1.304322488117321e+17, 1.304322488207945e+17, 1.30432248829857e+17, 1.304322488389196e+17, 1.304322488479821e+17, 1.304322488570445e+17, 1.30432248866107e+17, 1.304322488751694e+17, 1.304322488842319e+17, 1.304322488932945e+17, 1.30432248902357e+17, 1.304322489112632e+17, 1.304322489203258e+17, 1.304322489293883e+17, 1.304322489384508e+17, 1.304322489475132e+17, 1.304322489564195e+17, 1.304322489656383e+17, 1.304322489747008e+17, 1.304322489837632e+17, 1.304322489928257e+17, 1.304322490018883e+17, 1.304322490107945e+17, 1.30432249019857e+17, 1.304322490289194e+17, 1.30432249037982e+17, 1.304322490470445e+17, 1.30432249056107e+17, 1.304322490651695e+17, 1.304322490740758e+17, 1.304322490832945e+17, 1.30432249092357e+17, 1.304322491012632e+17, 1.304322491103258e+17, 1.304322491193882e+17, 1.304322491284507e+17, 1.304322491375132e+17, 1.304322491465757e+17, 1.304322491556383e+17, 1.304322491647008e+17, 1.304322491737633e+17, 1.304322491828257e+17, 1.30432249191732e+17, 1.304322492007945e+17, 1.30432249209857e+17, 1.304322492189196e+17, 1.30432249227982e+17, 1.304322492370445e+17, 1.30432249246107e+17, 1.304322492551695e+17, 1.304322492642321e+17, 1.304322492732945e+17, 1.30432249282357e+17, 1.304322492912632e+17, 1.304322493003256e+17, 1.304322493093883e+17, 1.304322493184507e+17, 1.304322493275132e+17, 1.304322493364196e+17, 1.30432249345482e+17, 1.304322493545445e+17, 1.304322493637633e+17, 1.304322493726694e+17, 1.30432249381732e+17, 1.304322493907945e+17, 1.30432249399857e+17, 1.304322494089196e+17, 1.304322494179821e+17, 1.304322494270445e+17, 1.30432249436107e+17, 1.304322494451695e+17, 1.304322494542321e+17, 1.304322494632945e+17, 1.30432249472357e+17, 1.304322494814194e+17, 1.304322494904819e+17, 1.304322494995444e+17, 1.304322495084508e+17, 1.304322495175133e+17, 1.304322495265757e+17, 1.304322495356383e+17, 1.304322495447007e+17, 1.304322495537632e+17, 1.304322495628257e+17, 1.30432249571732e+17, 1.304322495807945e+17, 1.304322495900133e+17, 1.304322495990757e+17, 1.304322496079821e+17, 1.304322496170445e+17, 1.30432249626107e+17, 1.304322496351695e+17, 1.304322496442319e+17, 1.304322496531383e+17, 1.30432249662357e+17, 1.304322496714195e+17, 1.30432249680482e+17, 1.304322496895444e+17, 1.304322496984508e+17, 1.304322497075132e+17, 1.304322497165757e+17, 1.304322497256381e+17, 1.304322497347007e+17, 1.304322497437632e+17, 1.304322497526696e+17, 1.30432249761732e+17, 1.304322497707945e+17, 1.30432249779857e+17, 1.304322497889194e+17, 1.304322497978257e+17, 1.304322498068882e+17, 1.304322498159507e+17, 1.304322498250132e+17, 1.304322498340758e+17, 1.304322498431383e+17, 1.304322498522008e+17, 1.304322498614195e+17, 1.304322498703258e+17, 1.304322498795446e+17, 1.30432249888607e+17, 1.304322498976695e+17, 1.304322499065757e+17, 1.304322499156383e+17, 1.304322499247008e+17, 1.304322499337632e+17, 1.304322499428257e+17, 1.304322499518883e+17, 1.304322499611071e+17, 1.304322499700133e+17, 1.30432249979232e+17, 1.304322499882945e+17, 1.304322499973571e+17, 1.304322500064195e+17, 1.304322500153257e+17, 1.304322500243882e+17, 1.304322500334508e+17, 1.304322500425133e+17, 1.304322500515757e+17, 1.304322500606383e+17, 1.304322500697007e+17, 1.304322500787633e+17, 1.304322500878258e+17, 1.304322500968882e+17, 1.304322501057944e+17, 1.30432250114857e+17, 1.304322501239195e+17, 1.30432250132982e+17, 1.304322501420445e+17, 1.304322501511071e+17, 1.304322501601695e+17, 1.304322501690757e+17, 1.304322501781382e+17, 1.304322501872008e+17, 1.304322501962633e+17, 1.304322502053258e+17, 1.304322502143884e+17, 1.304322502234508e+17, 1.304322502325133e+17, 1.304322502415758e+17, 1.304322502506382e+17, 1.304322502597007e+17, 1.304322502687633e+17, 1.304322502778257e+17, 1.304322502868882e+17, 1.304322502959507e+17, 1.304322503050132e+17, 1.304322503139195e+17, 1.30432250322982e+17, 1.304322503320445e+17, 1.304322503411069e+17, 1.304322503501695e+17, 1.30432250359232e+17, 1.304322503681382e+17, 1.304322503773571e+17, 1.304322503862633e+17, 1.30432250395482e+17, 1.304322504045445e+17, 1.304322504134508e+17, 1.304322504225133e+17, 1.304322504315757e+17, 1.304322504406382e+17, 1.304322504497007e+17, 1.304322504587633e+17, 1.304322504678257e+17, 1.304322504768882e+17, 1.304322504859507e+17, 1.304322504950132e+17, 1.304322505040758e+17, 1.304322505129819e+17, 1.304322505220444e+17, 1.304322505311069e+17, 1.304322505401695e+17, 1.30432250549232e+17, 1.304322505582945e+17, 1.304322505673571e+17, 1.304322505764196e+17, 1.304322505854821e+17, 1.304322505945445e+17, 1.30432250603607e+17, 1.304322506125133e+17, 1.304322506215757e+17, 1.304322506306383e+17, 1.304322506397007e+17, 1.304322506487633e+17, 1.304322506576695e+17, 1.30432250666732e+17, 1.304322506759508e+17, 1.304322506850132e+17, 1.304322506940756e+17, 1.30432250702982e+17, 1.304322507120444e+17, 1.304322507211069e+17, 1.304322507301695e+17, 1.30432250739232e+17, 1.304322507481382e+17, 1.304322507572006e+17, 1.304322507662632e+17, 1.304322507753257e+17, 1.304322507843882e+17, 1.304322507934508e+17, 1.30432250802357e+17, 1.304322508114195e+17, 1.30432250820482e+17, 1.304322508295444e+17, 1.30432250838607e+17, 1.304322508476695e+17, 1.30432250856732e+17, 1.304322508657944e+17, 1.304322508748571e+17, 1.304322508839195e+17, 1.304322508928257e+17, 1.304322509018883e+17, 1.304322509109508e+17, 1.304322509200132e+17, 1.304322509290757e+17, 1.304322509381382e+17, 1.304322509472008e+17, 1.304322509562633e+17, 1.304322509653257e+17, 1.304322509742321e+17, 1.304322509834508e+17, 1.304322509925133e+17, 1.304322510015758e+17, 1.304322510104819e+17, 1.304322510197007e+17, 1.30432251028607e+17, 1.304322510376695e+17, 1.30432251046732e+17, 1.304322510557946e+17, 1.304322510648571e+17, 1.304322510739196e+17, 1.30432251082982e+17, 1.304322510920445e+17, 1.304322511011069e+17, 1.304322511101695e+17, 1.30432251119232e+17, 1.304322511282944e+17, 1.304322511373569e+17, 1.304322511464195e+17, 1.30432251155482e+17, 1.304322511645445e+17, 1.30432251173607e+17, 1.304322511826696e+17, 1.304322511915757e+17, 1.304322512006382e+17, 1.304322512097007e+17, 1.304322512187633e+17, 1.304322512278258e+17, 1.304322512368883e+17, 1.304322512457946e+17, 1.30432251254857e+17, 1.304322512639195e+17, 1.30432251272982e+17, 1.304322512820444e+17, 1.304322512911069e+17, 1.304322513000133e+17, 1.304322513090758e+17, 1.304322513181384e+17, 1.304322513272008e+17, 1.304322513362633e+17, 1.304322513453257e+17, 1.304322513543882e+17, 1.304322513634508e+17, 1.304322513725133e+17, 1.304322513815757e+17, 1.304322513906382e+17, 1.304322513995444e+17, 1.30432251408607e+17, 1.304322514176695e+17, 1.304322514267319e+17, 1.304322514357944e+17, 1.30432251444857e+17, 1.304322514539195e+17, 1.30432251462982e+17, 1.304322514720445e+17, 1.304322514811071e+17, 1.304322514901696e+17, 1.30432251499232e+17, 1.304322515081382e+17, 1.304322515172008e+17, 1.304322515262633e+17, 1.304322515353257e+17, 1.304322515443882e+17, 1.304322515534508e+17, 1.304322515625133e+17, 1.304322515715757e+17, 1.304322515806383e+17, 1.304322515895444e+17, 1.30432251598607e+17, 1.304322516076695e+17, 1.30432251616732e+17, 1.304322516256383e+17, 1.304322516347008e+17, 1.304322516437633e+17, 1.30432251652982e+17, 1.304322516618883e+17, 1.304322516709507e+17, 1.304322516801696e+17, 1.304322516890757e+17, 1.304322516981382e+17, 1.304322517072008e+17, 1.304322517162633e+17, 1.304322517253257e+17, 1.304322517342321e+17, 1.304322517432945e+17, 1.304322517525133e+17, 1.304322517614195e+17, 1.304322517706382e+17, 1.304322517797007e+17, 1.304322517887631e+17, 1.304322517976695e+17, 1.30432251806732e+17, 1.304322518157944e+17, 1.30432251824857e+17, 1.304322518339195e+17, 1.30432251842982e+17, 1.304322518520445e+17, 1.304322518609507e+17, 1.304322518701695e+17, 1.30432251879232e+17, 1.304322518882945e+17, 1.304322518972008e+17, 1.304322519062633e+17, 1.304322519153258e+17, 1.304322519243884e+17, 1.304322519332945e+17, 1.30432251942357e+17, 1.304322519514195e+17, 1.30432251960482e+17, 1.304322519695444e+17, 1.304322519787633e+17, 1.304322519878257e+17, 1.30432251996732e+17, 1.304322520057946e+17, 1.30432252014857e+17, 1.304322520239195e+17, 1.304322520329819e+17, 1.304322520420444e+17, 1.304322520509508e+17, 1.304322520600133e+17, 1.304322520690757e+17, 1.304322520782945e+17, 1.304322520872008e+17, 1.304322520962633e+17, 1.304322521053257e+17, 1.304322521143882e+17, 1.304322521234508e+17, 1.304322521325133e+17, 1.304322521414195e+17, 1.304322521506382e+17, 1.304322521597007e+17, 1.304322521687633e+17, 1.304322521778258e+17, 1.30432252186732e+17, 1.304322521957944e+17, 1.30432252204857e+17, 1.304322522139195e+17, 1.30432252222982e+17, 1.304322522318883e+17, 1.304322522411069e+17, 1.304322522501695e+17, 1.30432252259232e+17, 1.304322522682945e+17, 1.304322522773571e+17, 1.304322522864195e+17, 1.30432252295482e+17, 1.304322523045445e+17, 1.30432252313607e+17, 1.304322523226694e+17, 1.30432252331732e+17, 1.304322523406383e+17, 1.304322523497009e+17, 1.304322523587633e+17, 1.304322523679821e+17, 1.304322523768882e+17, 1.304322523859507e+17, 1.304322523951695e+17, 1.304322524040756e+17, 1.304322524131382e+17, 1.304322524222007e+17, 1.304322524312632e+17, 1.304322524403258e+17, 1.30432252449232e+17, 1.304322524582945e+17, 1.304322524675133e+17, 1.304322524765757e+17, 1.30432252485482e+17, 1.304322524947007e+17, 1.30432252503607e+17, 1.304322525126696e+17, 1.304322525217321e+17, 1.304322525307945e+17, 1.30432252539857e+17, 1.304322525487633e+17, 1.304322525578257e+17, 1.304322525668882e+17, 1.304322525759507e+17, 1.304322525850132e+17, 1.304322525939196e+17, 1.30432252602982e+17, 1.304322526120445e+17, 1.304322526211069e+17, 1.304322526301695e+17, 1.30432252639232e+17, 1.304322526482944e+17, 1.304322526572008e+17, 1.304322526664195e+17, 1.304322526753257e+17, 1.304322526843884e+17, 1.304322526934508e+17, 1.304322527025133e+17, 1.304322527115757e+17, 1.304322527206382e+17, 1.304322527297007e+17, 1.304322527387633e+17, 1.304322527478258e+17, 1.304322527568883e+17, 1.304322527659508e+17, 1.304322527750132e+17, 1.304322527839195e+17, 1.30432252792982e+17, 1.304322528020444e+17, 1.304322528111069e+17, 1.304322528201695e+17, 1.30432252829232e+17, 1.304322528382945e+17, 1.304322528473571e+17, 1.304322528564195e+17, 1.30432252865482e+17, 1.304322528745445e+17, 1.304322528834508e+17, 1.304322528925133e+17, 1.304322529015757e+17, 1.304322529106382e+17, 1.304322529197007e+17, 1.304322529286071e+17, 1.304322529376695e+17, 1.30432252946732e+17, 1.304322529557944e+17, 1.30432252964857e+17, 1.304322529737632e+17, 1.304322529828257e+17, 1.304322529918883e+17, 1.304322530009508e+17, 1.304322530100133e+17, 1.304322530190757e+17, 1.304322530281382e+17, 1.304322530372008e+17, 1.304322530464195e+17, 1.30432253055482e+17, 1.304322530645444e+17, 1.304322530736069e+17, 1.304322530826694e+17, 1.304322530915757e+17, 1.304322531006382e+17, 1.304322531097007e+17, 1.304322531187633e+17, 1.304322531278258e+17, 1.304322531368882e+17, 1.304322531459507e+17, 1.304322531550132e+17, 1.304322531640758e+17, 1.30432253172982e+17, 1.304322531820445e+17, 1.304322531911071e+17, 1.304322532001696e+17, 1.30432253209232e+17, 1.304322532182945e+17, 1.304322532272008e+17, 1.304322532362633e+17, 1.30432253245482e+17, 1.304322532545445e+17, 1.30432253263607e+17, 1.304322532726694e+17, 1.30432253281732e+17, 1.304322532906382e+17, 1.304322532997007e+17, 1.304322533089196e+17, 1.304322533178257e+17, 1.304322533268882e+17, 1.304322533359507e+17, 1.304322533450132e+17, 1.304322533540758e+17, 1.304322533631383e+17, 1.304322533722008e+17, 1.304322533812634e+17, 1.304322533901695e+17, 1.30432253399232e+17, 1.304322534082945e+17, 1.304322534173571e+17, 1.304322534264195e+17, 1.30432253435482e+17, 1.304322534443884e+17, 1.304322534534508e+17, 1.304322534626696e+17, 1.304322534717321e+17, 1.304322534807945e+17, 1.304322534897007e+17, 1.304322534987633e+17, 1.304322535078257e+17, 1.304322535168882e+17, 1.304322535259507e+17, 1.304322535350132e+17, 1.304322535440758e+17, 1.304322535531383e+17, 1.304322535622008e+17, 1.304322535712632e+17, 1.304322535803258e+17, 1.30432253589232e+17, 1.304322535982945e+17, 1.304322536073571e+17, 1.304322536164196e+17, 1.304322536254821e+17, 1.304322536345445e+17, 1.30432253643607e+17, 1.304322536526694e+17, 1.30432253661732e+17, 1.304322536707944e+17, 1.304322536797007e+17, 1.304322536887633e+17, 1.304322536978258e+17, 1.304322537068883e+17, 1.304322537159508e+17, 1.304322537250132e+17, 1.304322537340758e+17, 1.304322537431382e+17, 1.304322537522007e+17, 1.304322537612632e+17, 1.304322537703258e+17, 1.304322537793883e+17, 1.304322537882945e+17, 1.304322537973571e+17, 1.304322538064196e+17, 1.30432253815482e+17, 1.304322538245445e+17, 1.30432253833607e+17, 1.304322538426694e+17, 1.30432253851732e+17, 1.304322538607945e+17, 1.30432253869857e+17, 1.304322538789196e+17, 1.304322538878258e+17, 1.304322538968882e+17, 1.304322539059507e+17, 1.304322539150132e+17, 1.304322539240756e+17, 1.304322539331382e+17, 1.304322539422007e+17, 1.304322539512632e+17, 1.304322539603258e+17, 1.304322539693883e+17, 1.304322539784508e+17, 1.304322539875133e+17, 1.304322539964195e+17, 1.304322540056383e+17, 1.304322540145445e+17, 1.30432254023607e+17, 1.304322540326696e+17, 1.304322540417321e+17, 1.304322540507945e+17, 1.30432254059857e+17, 1.304322540689196e+17, 1.304322540779821e+17, 1.304322540870445e+17, 1.304322540959507e+17, 1.304322541050132e+17, 1.304322541140758e+17, 1.304322541231383e+17, 1.304322541322007e+17, 1.304322541412632e+17, 1.304322541503258e+17, 1.30432254159232e+17, 1.304322541684507e+17, 1.304322541773569e+17, 1.304322541864195e+17, 1.30432254195482e+17, 1.304322542045445e+17, 1.30432254213607e+17, 1.304322542226696e+17, 1.304322542315757e+17, 1.304322542407945e+17, 1.30432254249857e+17, 1.304322542589194e+17, 1.30432254267982e+17, 1.304322542770445e+17, 1.304322542859508e+17, 1.304322542950132e+17, 1.304322543040758e+17, 1.304322543131383e+17, 1.304322543222008e+17, 1.304322543312632e+17, 1.304322543401695e+17, 1.30432254349232e+17, 1.304322543584507e+17, 1.304322543675132e+17, 1.304322543764195e+17, 1.30432254385482e+17, 1.304322543945445e+17, 1.30432254403607e+17, 1.304322544126694e+17, 1.30432254421732e+17, 1.304322544306382e+17, 1.30432254439857e+17, 1.304322544487633e+17, 1.304322544578258e+17, 1.304322544670445e+17, 1.304322544759508e+17, 1.304322544850132e+17, 1.304322544940758e+17, 1.304322545031382e+17, 1.304322545122007e+17, 1.304322545212632e+17, 1.304322545303258e+17, 1.304322545393883e+17, 1.304322545484507e+17, 1.304322545575132e+17, 1.304322545665757e+17, 1.304322545756383e+17, 1.304322545845445e+17, 1.304322545936069e+17, 1.304322546026694e+17, 1.30432254611732e+17, 1.304322546207945e+17, 1.30432254629857e+17, 1.304322546389196e+17, 1.304322546479821e+17, 1.304322546570445e+17, 1.30432254666107e+17, 1.304322546750132e+17, 1.304322546840758e+17, 1.304322546931383e+17, 1.304322547022007e+17, 1.304322547112632e+17, 1.304322547203258e+17, 1.304322547293883e+17, 1.304322547384508e+17, 1.304322547475133e+17, 1.304322547565757e+17, 1.304322547656383e+17, 1.304322547745444e+17, 1.30432254783607e+17, 1.304322547926694e+17, 1.30432254801732e+17, 1.304322548107945e+17, 1.304322548197007e+17, 1.304322548287633e+17, 1.304322548379821e+17, 1.304322548470445e+17, 1.30432254856107e+17, 1.304322548651695e+17, 1.304322548742319e+17, 1.304322548831383e+17, 1.304322548922008e+17, 1.304322549012634e+17, 1.304322549103258e+17, 1.304322549193883e+17, 1.304322549284508e+17, 1.304322549375132e+17, 1.304322549465756e+17, 1.304322549556383e+17, 1.304322549647007e+17, 1.304322549737632e+17, 1.304322549826696e+17, 1.304322549917321e+17, 1.304322550007945e+17, 1.30432255009857e+17, 1.304322550189194e+17, 1.30432255027982e+17, 1.304322550370445e+17, 1.30432255046107e+17, 1.304322550553257e+17, 1.304322550642321e+17, 1.304322550734508e+17, 1.304322550825133e+17, 1.304322550915757e+17, 1.304322551006382e+17, 1.304322551097007e+17, 1.304322551187633e+17, 1.304322551276695e+17, 1.304322551367319e+17, 1.304322551457944e+17, 1.30432255154857e+17, 1.304322551639195e+17, 1.30432255172982e+17, 1.304322551820445e+17, 1.304322551911071e+17, 1.304322552001696e+17, 1.30432255209232e+17, 1.304322552182945e+17, 1.304322552272008e+17, 1.304322552362633e+17, 1.304322552453257e+17, 1.304322552543882e+17, 1.304322552634508e+17, 1.304322552725133e+17, 1.304322552815758e+17, 1.304322552906383e+17, 1.304322552997007e+17, 1.304322553087633e+17, 1.304322553178257e+17, 1.304322553268882e+17, 1.304322553357944e+17, 1.30432255344857e+17, 1.304322553539195e+17, 1.30432255362982e+17, 1.304322553720445e+17, 1.304322553811071e+17, 1.304322553901695e+17, 1.30432255399232e+17, 1.304322554082944e+17, 1.304322554173569e+17, 1.304322554264195e+17, 1.30432255435482e+17, 1.304322554443884e+17, 1.304322554534508e+17, 1.304322554625133e+17, 1.30432255471732e+17, 1.304322554806382e+17, 1.30432255489857e+17, 1.304322554989196e+17, 1.304322555078257e+17, 1.304322555168882e+17, 1.304322555259507e+17, 1.304322555350132e+17, 1.304322555440758e+17, 1.304322555531383e+17, 1.304322555620444e+17, 1.304322555712634e+17, 1.304322555803258e+17, 1.304322555895444e+17, 1.304322555984507e+17, 1.304322556075132e+17, 1.304322556165757e+17, 1.304322556256383e+17, 1.304322556347008e+17, 1.304322556437632e+17, 1.304322556528257e+17, 1.30432255661732e+17, 1.304322556707945e+17, 1.304322556798569e+17, 1.304322556889194e+17, 1.304322556978257e+17, 1.304322557068883e+17, 1.304322557159507e+17, 1.304322557250132e+17, 1.304322557340758e+17, 1.304322557431383e+17, 1.304322557520444e+17, 1.304322557612632e+17, 1.304322557703258e+17, 1.30432255779232e+17, 1.304322557884508e+17, 1.304322557975132e+17, 1.304322558064196e+17, 1.304322558154821e+17, 1.304322558245445e+17, 1.30432255833607e+17, 1.304322558426694e+17, 1.30432255851732e+17, 1.304322558606383e+17, 1.30432255869857e+17, 1.304322558789194e+17, 1.304322558878258e+17, 1.304322558968883e+17, 1.304322559059507e+17, 1.304322559150132e+17, 1.304322559240756e+17, 1.30432255932982e+17, 1.304322559422007e+17, 1.304322559511071e+17, 1.304322559601695e+17, 1.304322559693883e+17, 1.304322559782945e+17, 1.304322559873571e+17, 1.304322559964195e+17, 1.30432256005482e+17, 1.304322560145445e+17, 1.30432256023607e+17, 1.304322560326696e+17, 1.30432256041732e+17, 1.304322560506383e+17, 1.304322560597009e+17, 1.304322560689196e+17, 1.304322560779821e+17, 1.304322560870445e+17, 1.304322560959507e+17, 1.304322561050132e+17, 1.304322561140756e+17, 1.304322561231382e+17, 1.304322561322007e+17, 1.304322561412632e+17, 1.304322561503258e+17, 1.304322561593883e+17, 1.304322561684508e+17, 1.304322561775132e+17, 1.304322561865757e+17, 1.30432256195482e+17, 1.304322562045445e+17, 1.30432256213607e+17, 1.304322562226696e+17, 1.304322562317321e+17, 1.304322562407945e+17, 1.30432256249857e+17, 1.304322562589196e+17, 1.30432256267982e+17, 1.304322562770445e+17, 1.30432256286107e+17, 1.304322562950132e+17, 1.304322563040758e+17, 1.304322563131383e+17, 1.304322563222008e+17, 1.304322563312632e+17, 1.304322563401695e+17, 1.30432256349232e+17, 1.304322563582944e+17, 1.304322563675132e+17, 1.304322563764195e+17, 1.304322563856383e+17, 1.304322563945445e+17, 1.30432256403607e+17, 1.304322564126696e+17, 1.30432256421732e+17, 1.304322564307945e+17, 1.30432256439857e+17, 1.304322564487633e+17, 1.304322564578258e+17, 1.304322564670445e+17, 1.30432256476107e+17, 1.304322564851695e+17, 1.304322564940758e+17, 1.304322565031383e+17, 1.304322565122007e+17, 1.304322565212632e+17, 1.304322565303256e+17, 1.304322565393882e+17, 1.304322565482945e+17, 1.304322565573571e+17, 1.304322565665757e+17, 1.304322565756383e+17, 1.304322565845445e+17, 1.304322565937633e+17, 1.304322566026694e+17, 1.30432256611732e+17, 1.304322566207945e+17, 1.30432256629857e+17, 1.304322566389196e+17, 1.304322566478258e+17, 1.304322566568883e+17, 1.30432256666107e+17, 1.304322566750132e+17, 1.304322566840756e+17, 1.304322566931382e+17, 1.304322567022007e+17, 1.304322567112632e+17, 1.304322567203258e+17, 1.30432256729232e+17, 1.304322567382945e+17, 1.304322567473571e+17, 1.304322567564195e+17, 1.304322567656383e+17, 1.304322567745444e+17, 1.304322567837632e+17, 1.304322567926694e+17, 1.30432256801732e+17, 1.304322568107945e+17, 1.30432256819857e+17, 1.304322568289196e+17, 1.304322568378258e+17, 1.304322568468882e+17, 1.304322568559507e+17, 1.304322568651695e+17, 1.304322568740758e+17, 1.304322568832945e+17, 1.304322568922008e+17, 1.304322569012632e+17, 1.304322569103258e+17, 1.304322569193883e+17, 1.304322569284508e+17, 1.304322569373569e+17, 1.304322569464195e+17, 1.30432256955482e+17, 1.304322569647007e+17, 1.304322569737632e+17, 1.30432256982982e+17, 1.304322569920444e+17, 1.304322570009508e+17, 1.304322570100133e+17, 1.304322570190757e+17, 1.304322570281384e+17, 1.304322570372008e+17, 1.304322570462633e+17, 1.304322570551695e+17, 1.304322570642321e+17, 1.304322570732945e+17, 1.304322570825132e+17, 1.304322570915757e+17, 1.304322571006382e+17, 1.304322571097007e+17, 1.30432257118607e+17, 1.304322571276695e+17, 1.30432257136732e+17, 1.304322571457944e+17, 1.30432257154857e+17, 1.304322571637632e+17, 1.304322571728257e+17, 1.304322571820445e+17, 1.304322571911071e+17, 1.304322572001695e+17, 1.30432257209232e+17, 1.304322572181382e+17, 1.304322572272008e+17, 1.304322572362632e+17, 1.304322572453257e+17, 1.304322572543882e+17, 1.304322572632945e+17, 1.30432257272357e+17, 1.304322572815757e+17, 1.304322572906382e+17, 1.304322572995444e+17, 1.304322573087633e+17, 1.304322573176695e+17, 1.304322573267319e+17, 1.304322573357944e+17, 1.30432257344857e+17, 1.304322573539195e+17, 1.30432257362982e+17, 1.304322573720445e+17, 1.304322573811071e+17, 1.304322573901696e+17, 1.304322573993883e+17, 1.304322574082945e+17, 1.304322574175133e+17, 1.304322574265757e+17, 1.304322574357946e+17, 1.304322574448571e+17, 1.304322574539196e+17, 1.30432257462982e+17, 1.304322574720444e+17, 1.304322574811069e+17, 1.304322574901695e+17, 1.30432257499232e+17, 1.304322575082944e+17, 1.304322575173569e+17, 1.304322575262633e+17, 1.30432257535482e+17, 1.304322575445445e+17, 1.304322575537633e+17, 1.304322575626696e+17, 1.304322575718883e+17, 1.304322575807945e+17, 1.30432257589857e+17, 1.304322575989194e+17, 1.30432257607982e+17, 1.304322576170445e+17, 1.304322576259508e+17, 1.304322576350132e+17, 1.304322576440758e+17, 1.304322576532945e+17, 1.304322576622007e+17, 1.304322576714195e+17, 1.304322576803256e+17, 1.304322576893882e+17, 1.304322576984507e+17, 1.304322577075132e+17, 1.304322577165757e+17, 1.304322577256383e+17, 1.304322577345445e+17, 1.30432257743607e+17, 1.304322577528259e+17, 1.304322577618883e+17, 1.304322577709508e+17, 1.304322577800132e+17, 1.304322577890757e+17, 1.304322577979821e+17, 1.304322578070445e+17, 1.30432257816107e+17, 1.304322578251695e+17, 1.304322578342321e+17, 1.304322578432945e+17, 1.30432257852357e+17, 1.304322578614194e+17, 1.304322578704819e+17, 1.304322578795444e+17, 1.30432257888607e+17, 1.304322578975132e+17, 1.304322579065757e+17, 1.304322579156383e+17, 1.304322579247008e+17, 1.304322579337632e+17, 1.304322579428257e+17, 1.304322579518883e+17, 1.304322579609508e+17, 1.304322579700133e+17, 1.304322579790757e+17, 1.304322579881382e+17, 1.304322579972008e+17, 1.304322580062633e+17, 1.304322580153257e+17, 1.304322580243882e+17, 1.304322580334508e+17, 1.304322580425133e+17, 1.304322580514195e+17, 1.30432258060482e+17, 1.304322580697007e+17, 1.30432258078607e+17, 1.304322580878258e+17, 1.304322580968883e+17, 1.304322581057946e+17, 1.304322581148571e+17, 1.304322581239195e+17, 1.30432258132982e+17, 1.304322581420444e+17, 1.304322581511069e+17, 1.304322581601695e+17, 1.30432258169232e+17, 1.304322581782945e+17, 1.304322581873571e+17, 1.304322581964195e+17, 1.304322582053257e+17, 1.304322582143882e+17, 1.304322582234508e+17, 1.304322582325132e+17, 1.304322582415757e+17, 1.304322582506382e+17, 1.304322582597007e+17, 1.304322582687633e+17, 1.304322582778258e+17, 1.304322582868883e+17, 1.304322582957944e+17, 1.30432258304857e+17, 1.304322583139195e+17, 1.30432258322982e+17, 1.304322583320445e+17, 1.304322583411071e+17, 1.304322583501695e+17, 1.304322583590758e+17, 1.304322583682945e+17, 1.304322583773571e+17, 1.304322583864196e+17, 1.30432258395482e+17, 1.304322584043882e+17, 1.304322584134508e+17, 1.304322584225133e+17, 1.304322584315757e+17, 1.304322584406382e+17, 1.304322584497007e+17, 1.304322584587633e+17, 1.304322584678258e+17, 1.304322584768882e+17, 1.304322584859507e+17, 1.304322584950132e+17, 1.304322585039195e+17, 1.30432258512982e+17, 1.304322585220445e+17, 1.304322585311071e+17, 1.304322585401696e+17, 1.30432258549232e+17, 1.304322585582945e+17, 1.304322585673569e+17, 1.304322585762633e+17, 1.30432258585482e+17, 1.304322585943882e+17, 1.304322586034508e+17, 1.304322586125133e+17, 1.304322586215758e+17, 1.304322586306383e+17, 1.304322586397007e+17, 1.304322586487633e+17, 1.304322586578257e+17, 1.304322586668882e+17, 1.304322586757944e+17, 1.30432258684857e+17, 1.304322586939195e+17, 1.30432258702982e+17, 1.304322587120445e+17, 1.304322587211069e+17, 1.304322587301695e+17, 1.30432258739232e+17, 1.304322587482945e+17, 1.304322587572008e+17, 1.304322587664195e+17, 1.30432258775482e+17, 1.304322587845445e+17, 1.30432258793607e+17, 1.304322588026696e+17, 1.304322588117321e+17, 1.304322588207945e+17, 1.30432258829857e+17, 1.304322588389194e+17, 1.30432258847982e+17, 1.304322588568882e+17, 1.304322588659507e+17, 1.304322588750132e+17, 1.304322588840758e+17, 1.304322588931383e+17, 1.304322589020444e+17, 1.304322589111069e+17, 1.304322589201695e+17, 1.30432258929232e+17, 1.304322589382945e+17, 1.304322589473571e+17, 1.304322589564196e+17, 1.304322589654821e+17, 1.304322589745445e+17, 1.304322589837632e+17, 1.304322589928257e+17, 1.30432259001732e+17, 1.304322590109508e+17, 1.304322590198569e+17, 1.304322590289194e+17, 1.30432259037982e+17, 1.304322590470445e+17, 1.30432259056107e+17, 1.304322590650132e+17, 1.304322590740758e+17, 1.304322590832946e+17, 1.30432259092357e+17, 1.304322591014195e+17, 1.304322591104819e+17, 1.304322591193883e+17, 1.304322591284508e+17, 1.304322591375133e+17, 1.304322591465757e+17, 1.304322591556383e+17, 1.304322591645445e+17, 1.30432259173607e+17, 1.304322591828257e+17, 1.30432259191732e+17, 1.304322592007945e+17, 1.304322592095444e+17, 1.304322592178257e+17, 1.304322592257944e+17, 1.304322592334508e+17, 1.304322592475132e+17, 1.304322592607945e+17, 1.304322592737632e+17, 1.30432259285482e+17, 1.30432259296107e+17, 1.304322593062633e+17, 1.304322593162633e+17, 1.304322593264196e+17, 1.304322593364195e+17, 1.304322593464195e+17, 1.304322593564195e+17, 1.304322593664196e+17, 1.304322593765757e+17, 1.304322593865757e+17, 1.30432259396107e+17, 1.30432259404857e+17, 1.304322594131383e+17, 1.304322594211071e+17, 1.30432259429232e+17, 1.304322594373571e+17, 1.304322594453258e+17, 1.304322594532946e+17, 1.304322594614195e+17, 1.304322594693882e+17, 1.304322594775133e+17, 1.304322594851694e+17, 1.30432259495482e+17, 1.304322595047007e+17, 1.304322595134508e+17, 1.304322595218883e+17, 1.304322595314194e+17, 1.304322595407945e+17, 1.304322595482944e+17, 1.304322595557944e+17, 1.304322595634508e+17, 1.304322595709507e+17, 1.304322595784508e+17, 1.304322595859507e+17, 1.30432259593607e+17, 1.304322596012632e+17, 1.304322596087633e+17, 1.304322596162633e+17, 1.304322596239195e+17, 1.304322596339195e+17, 1.304322596412632e+17, 1.30432259648607e+17, 1.30432259656107e+17, 1.30432259663607e+17, 1.304322596709508e+17, 1.304322596784507e+17, 1.304322596857944e+17, 1.304322596931383e+17, 1.304322597006382e+17, 1.30432259707982e+17, 1.304322597151695e+17, 1.304322597225133e+17, 1.304322597300132e+17, 1.304322597373569e+17, 1.304322597447007e+17, 1.304322597520445e+17, 1.304322597593883e+17, 1.30432259766732e+17, 1.304322597742321e+17, 1.304322597818883e+17, 1.30432259789232e+17, 1.304322597965757e+17, 1.304322598039195e+17, 1.304322598114195e+17, 1.30432259818607e+17, 1.30432259826107e+17, 1.30432259833607e+17, 1.304322598409508e+17, 1.304322598482945e+17, 1.304322598556383e+17, 1.304322598631382e+17, 1.304322598704819e+17, 1.304322598779821e+17, 1.304322598851695e+17, 1.304322598925133e+17, 1.304322599000133e+17, 1.304322599073571e+17, 1.304322599147008e+17, 1.304322599222008e+17, 1.304322599297007e+17, 1.304322599370445e+17, 1.304322599443882e+17, 1.304322599515757e+17, 1.304322599589196e+17, 1.304322599662632e+17, 1.304322599737632e+17, 1.304322599814195e+17, 1.304322599887633e+17, 1.30432259996107e+17, 1.304322600034508e+17, 1.304322600107945e+17, 1.304322600181382e+17, 1.30432260025482e+17, 1.30432260032982e+17, 1.304322600401695e+17, 1.304322600475132e+17, 1.30432260054857e+17, 1.30432260062357e+17, 1.30432260069857e+17, 1.304322600773571e+17, 1.30432260084857e+17, 1.304322600920444e+17, 1.304322600993882e+17, 1.304322601067319e+17, 1.304322601142321e+17, 1.304322601215758e+17, 1.304322601289196e+17, 1.304322601362633e+17, 1.30432260143607e+17, 1.304322601509508e+17, 1.304322601582945e+17, 1.304322601656383e+17, 1.30432260172982e+17, 1.30432260180482e+17, 1.304322601876695e+17, 1.304322601951695e+17, 1.304322602025133e+17, 1.30432260209857e+17, 1.304322602172008e+17, 1.304322602245444e+17, 1.304322602320445e+17, 1.304322602395444e+17, 1.304322602468883e+17, 1.304322602542321e+17, 1.30432260261732e+17, 1.304322602690757e+17, 1.304322602765757e+17, 1.304322602839195e+17, 1.304322602914195e+17, 1.304322602987633e+17, 1.30432260306107e+17, 1.304322603134508e+17, 1.304322603207945e+17, 1.304322603284507e+17, 1.304322603357944e+17, 1.304322603431383e+17, 1.30432260350482e+17, 1.304322603578258e+17, 1.304322603651695e+17, 1.30432260372357e+17, 1.30432260379857e+17, 1.304322603873569e+17, 1.304322603947007e+17, 1.304322604020444e+17, 1.304322604093883e+17, 1.30432260416732e+17, 1.304322604240758e+17, 1.30432260431732e+17, 1.304322604390757e+17, 1.304322604464195e+17, 1.304322604537633e+17, 1.304322604609507e+17, 1.304322604684508e+17, 1.304322604757946e+17, 1.304322604831383e+17, 1.304322604903258e+17, 1.304322604978258e+17, 1.304322605053257e+17, 1.304322605126696e+17, 1.304322605200133e+17, 1.304322605275132e+17, 1.30432260534857e+17, 1.304322605422007e+17, 1.304322605495444e+17, 1.304322605568882e+17, 1.304322605640756e+17, 1.304322605715758e+17, 1.304322605790757e+17, 1.304322605864196e+17, 1.304322605939195e+17, 1.304322606014195e+17, 1.304322606087633e+17, 1.30432260616107e+17, 1.304322606234508e+17, 1.304322606309508e+17, 1.304322606382944e+17, 1.30432260645482e+17, 1.304322606528257e+17, 1.304322606601695e+17, 1.304322606676695e+17, 1.304322606750132e+17, 1.304322606825133e+17, 1.304322606900132e+17, 1.304322606973571e+17, 1.304322607048571e+17, 1.30432260712357e+17, 1.304322607197007e+17, 1.304322607272008e+17, 1.304322607347008e+17, 1.304322607422007e+17, 1.304322607493883e+17, 1.30432260756732e+17, 1.304322607642321e+17, 1.30432260771732e+17, 1.304322607790757e+17, 1.304322607864195e+17, 1.304322607937632e+17, 1.304322608011069e+17, 1.304322608084507e+17, 1.304322608159508e+17, 1.304322608232945e+17, 1.304322608307945e+17, 1.304322608382945e+17, 1.304322608456383e+17, 1.30432260852982e+17, 1.304322608603258e+17, 1.304322608676695e+17, 1.304322608751695e+17, 1.304322608825133e+17, 1.30432260889857e+17, 1.304322608972008e+17, 1.304322609045445e+17, 1.304322609118883e+17, 1.30432260919232e+17, 1.304322609265757e+17, 1.304322609342319e+17, 1.304322609417321e+17, 1.304322609489196e+17, 1.304322609562633e+17, 1.30432260963607e+17, 1.304322609712632e+17, 1.30432260978607e+17, 1.304322609859508e+17, 1.304322609931382e+17, 1.30432261000482e+17, 1.304322610078258e+17, 1.304322610150132e+17, 1.30432261022357e+17, 1.304322610297009e+17, 1.304322610372008e+17, 1.304322610443884e+17, 1.304322610518883e+17, 1.30432261059232e+17, 1.304322610665756e+17, 1.304322610739195e+17, 1.304322610815758e+17, 1.304322610889196e+17, 1.304322610962633e+17, 1.304322611037632e+17, 1.304322611111071e+17, 1.30432261118607e+17, 1.30432261126107e+17, 1.30432261133607e+17, 1.304322611409508e+17, 1.304322611484507e+17, 1.304322611556383e+17, 1.30432261162982e+17, 1.304322611703258e+17, 1.304322611776695e+17, 1.304322611850132e+17, 1.30432261192357e+17, 1.30432261199857e+17, 1.304322612072008e+17, 1.304322612145445e+17, 1.304322612218883e+17, 1.30432261229232e+17, 1.30432261236732e+17, 1.304322612440758e+17, 1.304322612515757e+17, 1.304322612589196e+17, 1.30432261266107e+17, 1.304322612734508e+17, 1.304322612811069e+17, 1.304322612884508e+17, 1.304322612957946e+17, 1.304322613032945e+17, 1.304322613106382e+17, 1.304322613181382e+17, 1.304322613253257e+17, 1.304322613328257e+17, 1.304322613401695e+17, 1.304322613475132e+17, 1.304322613547008e+17, 1.304322613622007e+17, 1.304322613695444e+17, 1.304322613768882e+17, 1.304322613843882e+17, 1.30432261391732e+17, 1.304322613990758e+17, 1.304322614064196e+17, 1.304322614137633e+17, 1.304322614212632e+17, 1.30432261428607e+17, 1.30432261436107e+17, 1.304322614434508e+17, 1.304322614507945e+17, 1.304322614581382e+17, 1.30432261465482e+17, 1.304322614728257e+17, 1.304322614803258e+17, 1.304322614876695e+17, 1.30432261494857e+17, 1.304322615023571e+17, 1.304322615097009e+17, 1.304322615168883e+17, 1.304322615242321e+17, 1.304322615318883e+17, 1.30432261539232e+17, 1.304322615465757e+17, 1.304322615540758e+17, 1.304322615615757e+17, 1.304322615689196e+17, 1.304322615762633e+17, 1.304322615837633e+17, 1.304322615912632e+17, 1.304322615984508e+17, 1.304322616059507e+17, 1.304322616132945e+17, 1.304322616204819e+17, 1.30432261627982e+17, 1.304322616353257e+17, 1.304322616428257e+17, 1.304322616501695e+17, 1.304322616575132e+17, 1.304322616650132e+17, 1.304322616725133e+17, 1.304322616800133e+17, 1.304322616873571e+17, 1.304322616947008e+17, 1.304322617022008e+17, 1.304322617095444e+17, 1.30432261716732e+17, 1.304322617242321e+17, 1.304322617320445e+17, 1.304322617393883e+17, 1.30432261746732e+17, 1.304322617540758e+17, 1.304322617614195e+17, 1.304322617687633e+17, 1.30432261776107e+17, 1.30432261783607e+17, 1.304322617909508e+17, 1.304322617982945e+17, 1.304322618056383e+17, 1.304322618131383e+17, 1.304322618203258e+17, 1.304322618276695e+17, 1.304322618350132e+17, 1.304322618425133e+17, 1.30432261849857e+17, 1.304322618572008e+17, 1.304322618645445e+17, 1.304322618718883e+17, 1.304322618795444e+17, 1.304322618868883e+17, 1.304322618942321e+17, 1.30432261901732e+17, 1.304322619090757e+17, 1.304322619162633e+17, 1.30432261923607e+17, 1.304322619312632e+17, 1.30432261938607e+17, 1.30432261946107e+17, 1.304322619536069e+17, 1.304322619609508e+17, 1.304322619682945e+17, 1.304322619757944e+17, 1.304322619832945e+17, 1.304322619904819e+17, 1.30432261997982e+17, 1.304322620051694e+17, 1.304322620125132e+17, 1.30432262019857e+17, 1.304322620270445e+17, 1.304322620345445e+17, 1.304322620418883e+17, 1.304322620490757e+17, 1.304322620564196e+17, 1.304322620639195e+17, 1.304322620712632e+17, 1.30432262078607e+17, 1.30432262086107e+17, 1.304322620934508e+17, 1.304322621006382e+17, 1.304322621079821e+17, 1.304322621153258e+17, 1.304322621228257e+17, 1.304322621303256e+17, 1.304322621378258e+17, 1.304322621451695e+17, 1.304322621526696e+17, 1.30432262159857e+17, 1.304322621672008e+17, 1.304322621745445e+17, 1.304322621818883e+17, 1.30432262189232e+17, 1.304322621964195e+17, 1.304322622037632e+17, 1.304322622111069e+17, 1.304322622184507e+17, 1.304322622259508e+17, 1.304322622331383e+17, 1.304322622406383e+17, 1.304322622479821e+17, 1.304322622553257e+17, 1.304322622625133e+17, 1.30432262269857e+17, 1.304322622773569e+17, 1.304322622847007e+17, 1.304322622918883e+17, 1.30432262299232e+17, 1.304322623065757e+17, 1.304322623139195e+17, 1.304322623212634e+17, 1.304322623286071e+17, 1.30432262336107e+17, 1.304322623436069e+17, 1.304322623509508e+17, 1.304322623581382e+17, 1.304322623656383e+17, 1.304322623731383e+17, 1.304322623806382e+17, 1.304322623881382e+17, 1.30432262395482e+17, 1.304322624028257e+17, 1.304322624101695e+17, 1.304322624175132e+17, 1.30432262424857e+17, 1.304322624322007e+17, 1.304322624397007e+17, 1.30432262447982e+17, 1.304322624553257e+17, 1.304322624626694e+17, 1.304322624701696e+17, 1.304322624775133e+17, 1.304322624850132e+17, 1.304322624922008e+17, 1.304322624997007e+17, 1.304322625070445e+17, 1.304322625143882e+17, 1.304322625218883e+17, 1.30432262529232e+17, 1.304322625365757e+17, 1.304322625440756e+17, 1.304322625515758e+17, 1.304322625587633e+17, 1.30432262566107e+17, 1.30432262573607e+17, 1.304322625812634e+17, 1.304322625886071e+17, 1.304322625959508e+17, 1.304322626034508e+17, 1.304322626107945e+17, 1.304322626181382e+17, 1.30432262625482e+17, 1.30432262632982e+17, 1.304322626403258e+17, 1.304322626475133e+17, 1.304322626550132e+17, 1.30432262662357e+17, 1.304322626697007e+17, 1.304322626772008e+17, 1.304322626847008e+17, 1.304322626922007e+17, 1.304322626993883e+17, 1.30432262706732e+17, 1.304322627140756e+17, 1.304322627214194e+17, 1.304322627287633e+17, 1.304322627362633e+17, 1.30432262743607e+17, 1.304322627511069e+17, 1.304322627584507e+17, 1.304322627656383e+17, 1.30432262772982e+17, 1.304322627803258e+17, 1.304322627876695e+17, 1.304322627950132e+17, 1.30432262802357e+17, 1.304322628097009e+17, 1.304322628170445e+17, 1.304322628243884e+17, 1.304322628318883e+17, 1.304322628393883e+17, 1.304322628465756e+17, 1.304322628540758e+17, 1.304322628615758e+17, 1.304322628689196e+17, 1.304322628762633e+17, 1.304322628839195e+17, 1.304322628912632e+17, 1.30432262898607e+17, 1.30432262906107e+17, 1.304322629134508e+17, 1.304322629207945e+17, 1.304322629284507e+17, 1.304322629357944e+17, 1.304322629431382e+17, 1.304322629506383e+17, 1.304322629579821e+17, 1.304322629653258e+17, 1.304322629726696e+17, 1.304322629800133e+17, 1.304322629873571e+17, 1.304322629947008e+17, 1.304322630020444e+17, 1.304322630097007e+17, 1.304322630170445e+17, 1.304322630245445e+17, 1.304322630322007e+17, 1.304322630395444e+17, 1.304322630468882e+17, 1.304322630543882e+17, 1.30432263061732e+17, 1.304322630690758e+17, 1.304322630764196e+17, 1.304322630839195e+17, 1.304322630911071e+17, 1.304322630984508e+17, 1.304322631057946e+17, 1.304322631132945e+17, 1.304322631206382e+17, 1.304322631281382e+17, 1.304322631356383e+17, 1.30432263142982e+17, 1.304322631503258e+17, 1.304322631576695e+17, 1.304322631650132e+17, 1.30432263172357e+17, 1.30432263179857e+17, 1.304322631872008e+17, 1.304322631945445e+17, 1.304322632018883e+17, 1.30432263209232e+17, 1.304322632164195e+17, 1.304322632237632e+17, 1.304322632311069e+17, 1.30432263238607e+17, 1.304322632459507e+17, 1.304322632532945e+17, 1.304322632607945e+17, 1.30432263267982e+17, 1.304322632753257e+17, 1.304322632828257e+17, 1.304322632901695e+17, 1.304322632973569e+17, 1.304322633047007e+17, 1.304322633122008e+17, 1.304322633193883e+17, 1.30432263326732e+17, 1.304322633342321e+17, 1.304322633415757e+17, 1.304322633490757e+17, 1.304322633564196e+17, 1.304322633637633e+17, 1.304322633712632e+17, 1.30432263378607e+17, 1.30432263386107e+17, 1.304322633934508e+17, 1.304322634009508e+17, 1.304322634082945e+17, 1.304322634157944e+17, 1.304322634231382e+17, 1.304322634306383e+17, 1.304322634379821e+17, 1.304322634453258e+17, 1.304322634528257e+17, 1.304322634601695e+17, 1.304322634675132e+17, 1.304322634751695e+17, 1.304322634825133e+17, 1.30432263489857e+17, 1.304322634972008e+17, 1.304322635045445e+17, 1.304322635118883e+17, 1.30432263519232e+17, 1.304322635265757e+17, 1.304322635340758e+17, 1.304322635415757e+17, 1.304322635489194e+17, 1.304322635562633e+17, 1.30432263563607e+17, 1.304322635709508e+17, 1.304322635784508e+17, 1.304322635859507e+17, 1.304322635931383e+17, 1.304322636006383e+17, 1.304322636081382e+17, 1.304322636153257e+17, 1.304322636225133e+17, 1.304322636300133e+17, 1.304322636375132e+17, 1.304322636447007e+17, 1.304322636520444e+17, 1.304322636593882e+17, 1.304322636667319e+17, 1.304322636740758e+17, 1.304322636815758e+17, 1.304322636890757e+17, 1.304322636964195e+17, 1.30432263703607e+17, 1.304322637111069e+17, 1.30432263718607e+17, 1.304322637259507e+17, 1.304322637342319e+17, 1.30432263741732e+17, 1.304322637490757e+17, 1.304322637564195e+17, 1.304322637637632e+17, 1.304322637712632e+17, 1.304322637784507e+17, 1.304322637859508e+17, 1.304322637931382e+17, 1.30432263800482e+17, 1.304322638079821e+17, 1.304322638153257e+17, 1.304322638226696e+17, 1.304322638300133e+17, 1.304322638376695e+17, 1.304322638448571e+17, 1.304322638520444e+17, 1.304322638595444e+17, 1.30432263866732e+17, 1.304322638742321e+17, 1.30432263881732e+17, 1.30432263889232e+17, 1.304322638965757e+17, 1.304322639039195e+17, 1.304322639115757e+17, 1.304322639189196e+17, 1.304322639262633e+17, 1.304322639337633e+17, 1.304322639412632e+17, 1.30432263948607e+17, 1.304322639559507e+17, 1.304322639632945e+17, 1.304322639706383e+17, 1.304322639779821e+17, 1.30432263985482e+17, 1.304322639928257e+17, 1.304322640001695e+17, 1.304322640075132e+17, 1.30432264014857e+17, 1.304322640220444e+17, 1.304322640293882e+17, 1.304322640367319e+17, 1.304322640440758e+17, 1.30432264051732e+17, 1.304322640590757e+17, 1.304322640664195e+17, 1.304322640737632e+17, 1.304322640811069e+17, 1.30432264088607e+17, 1.304322640959507e+17, 1.304322641032945e+17, 1.304322641106382e+17, 1.304322641181382e+17, 1.30432264125482e+17, 1.30432264132982e+17, 1.304322641403258e+17, 1.304322641476695e+17, 1.304322641550132e+17, 1.30432264162357e+17, 1.304322641697007e+17, 1.304322641770445e+17, 1.304322641845445e+17, 1.304322641918883e+17, 1.30432264199232e+17, 1.304322642065757e+17, 1.304322642139195e+17, 1.304322642212632e+17, 1.30432264228607e+17, 1.30432264236107e+17, 1.304322642434508e+17, 1.304322642507945e+17, 1.304322642581382e+17, 1.30432264265482e+17, 1.304322642728257e+17, 1.304322642801695e+17, 1.304322642875132e+17, 1.30432264294857e+17, 1.304322643022007e+17, 1.304322643097007e+17, 1.304322643170445e+17, 1.304322643243882e+17, 1.304322643320445e+17, 1.304322643393883e+17, 1.30432264346732e+17, 1.304322643542319e+17, 1.304322643626694e+17, 1.304322643700132e+17, 1.304322643772008e+17, 1.30432264384857e+17, 1.304322643922007e+17, 1.304322643993882e+17, 1.30432264406732e+17, 1.304322644140758e+17, 1.304322644215758e+17, 1.304322644289196e+17, 1.304322644364195e+17, 1.304322644437632e+17, 1.304322644511069e+17, 1.304322644584508e+17, 1.304322644657946e+17, 1.304322644731383e+17, 1.30432264480482e+17, 1.30432264487982e+17, 1.304322644953257e+17, 1.304322645028259e+17, 1.304322645100132e+17, 1.304322645173571e+17, 1.304322645248571e+17, 1.304322645322008e+17, 1.304322645395444e+17, 1.304322645468882e+17, 1.304322645542319e+17, 1.304322645617321e+17, 1.304322645690757e+17, 1.30432264576732e+17, 1.304322645840756e+17, 1.30432264591732e+17, 1.304322645989196e+17, 1.304322646064195e+17, 1.30432264613607e+17, 1.304322646209508e+17, 1.304322646286071e+17, 1.30432264636107e+17, 1.304322646432945e+17, 1.304322646506383e+17, 1.304322646579821e+17, 1.304322646653257e+17, 1.304322646726694e+17, 1.304322646801695e+17, 1.304322646876695e+17, 1.304322646950132e+17, 1.30432264702357e+17, 1.304322647097007e+17, 1.304322647168882e+17, 1.304322647242319e+17, 1.30432264731732e+17, 1.304322647390757e+17, 1.304322647464196e+17, 1.304322647537633e+17, 1.304322647611071e+17, 1.304322647684508e+17, 1.304322647756383e+17, 1.304322647832945e+17, 1.304322647906382e+17, 1.30432264797982e+17, 1.304322648053258e+17, 1.304322648126696e+17, 1.304322648200133e+17, 1.304322648276695e+17, 1.304322648351695e+17, 1.304322648425133e+17, 1.304322648500132e+17, 1.304322648573569e+17, 1.304322648647007e+17, 1.304322648720444e+17, 1.30432264879232e+17, 1.30432264886732e+17, 1.304322648940758e+17, 1.30432264901732e+17, 1.304322649090757e+17, 1.304322649162633e+17, 1.30432264923607e+17, 1.304322649309508e+17, 1.30432264938607e+17, 1.304322649457944e+17, 1.304322649531383e+17, 1.30432264960482e+17, 1.304322649678257e+17, 1.304322649751695e+17, 1.304322649825132e+17, 1.304322649900133e+17, 1.304322649975133e+17, 1.30432265004857e+17, 1.304322650122007e+17, 1.304322650195444e+17, 1.304322650268882e+17, 1.304322650343884e+17, 1.304322650420444e+17, 1.304322650493883e+17, 1.304322650565757e+17, 1.304322650640758e+17, 1.304322650715757e+17, 1.304322650789196e+17, 1.304322650864195e+17, 1.304322650937632e+17, 1.304322651011069e+17, 1.304322651084508e+17, 1.304322651157946e+17, 1.304322651232945e+17, 1.304322651306382e+17, 1.304322651382945e+17, 1.304322651456383e+17, 1.30432265152982e+17, 1.304322651603258e+17, 1.304322651676695e+17, 1.304322651751695e+17, 1.304322651825133e+17, 1.304322651900133e+17, 1.304322651973571e+17, 1.304322652047008e+17, 1.304322652120444e+17, 1.304322652193882e+17, 1.304322652267319e+17, 1.304322652342321e+17, 1.304322652420444e+17, 1.304322652493883e+17, 1.30432265256732e+17, 1.304322652640758e+17, 1.304322652714195e+17, 1.304322652787633e+17, 1.30432265286107e+17, 1.304322652937633e+17, 1.304322653011071e+17, 1.304322653084508e+17, 1.304322653156383e+17, 1.304322653231383e+17, 1.304322653303258e+17, 1.304322653376695e+17, 1.304322653450132e+17, 1.304322653525132e+17, 1.304322653598569e+17, 1.304322653672008e+17, 1.304322653745445e+17, 1.304322653822007e+17, 1.304322653895444e+17, 1.304322653968882e+17, 1.304322654043882e+17, 1.304322654118883e+17, 1.30432265419232e+17, 1.304322654265757e+17, 1.304322654339195e+17, 1.304322654415757e+17, 1.304322654487633e+17, 1.304322654562633e+17, 1.304322654634508e+17, 1.304322654709507e+17, 1.304322654784508e+17, 1.304322654859507e+17, 1.304322654932945e+17, 1.30432265500482e+17, 1.304322655078258e+17, 1.304322655151695e+17, 1.30432265522357e+17, 1.304322655297007e+17, 1.304322655370445e+17, 1.304322655445445e+17, 1.304322655518883e+17, 1.304322655593883e+17, 1.304322655665757e+17, 1.304322655739196e+17, 1.304322655812634e+17, 1.30432265588607e+17, 1.30432265596107e+17, 1.30432265603607e+17, 1.304322656109508e+17, 1.304322656182945e+17, 1.304322656256383e+17, 1.30432265632982e+17, 1.304322656403258e+17, 1.304322656476695e+17, 1.304322656550132e+17, 1.304322656625133e+17, 1.30432265669857e+17, 1.304322656772008e+17, 1.304322656845445e+17, 1.304322656922007e+17, 1.304322656995444e+17, 1.304322657068883e+17, 1.304322657142321e+17, 1.30432265721732e+17, 1.304322657290757e+17, 1.304322657364195e+17, 1.304322657439195e+17, 1.304322657512632e+17, 1.304322657584507e+17, 1.304322657659507e+17, 1.304322657732945e+17, 1.30432265780482e+17, 1.30432265787982e+17, 1.304322657953257e+17, 1.304322658028257e+17, 1.304322658101696e+17, 1.304322658175133e+17, 1.304322658250132e+17, 1.30432265832357e+17, 1.30432265839857e+17, 1.304322658472008e+17, 1.304322658545445e+17, 1.304322658618883e+17, 1.30432265869232e+17, 1.304322658765757e+17, 1.304322658840758e+17, 1.304322658915758e+17, 1.304322658987633e+17, 1.304322659062633e+17, 1.30432265913607e+17, 1.304322659209508e+17, 1.304322659284507e+17, 1.304322659359508e+17, 1.304322659432946e+17, 1.30432265950482e+17, 1.304322659578258e+17, 1.304322659653257e+17, 1.304322659725133e+17, 1.30432265979857e+17, 1.304322659873569e+17, 1.304322659947007e+17, 1.304322660020445e+17, 1.304322660093883e+17, 1.30432266016732e+17, 1.304322660243882e+17, 1.30432266031732e+17, 1.304322660392321e+17, 1.304322660465757e+17, 1.304322660539195e+17, 1.304322660612632e+17, 1.304322660687633e+17, 1.30432266076107e+17, 1.304322660834508e+17, 1.304322660911071e+17, 1.304322660984508e+17, 1.304322661057944e+17, 1.304322661132945e+17, 1.304322661204819e+17, 1.304322661278258e+17, 1.304322661351695e+17, 1.304322661426694e+17, 1.304322661500132e+17, 1.304322661573569e+17, 1.304322661647007e+17, 1.304322661720444e+17, 1.304322661795446e+17, 1.304322661868883e+17, 1.304322661943882e+17, 1.304322662018883e+17, 1.30432266209232e+17, 1.304322662164195e+17, 1.304322662239195e+17, 1.304322662312632e+17, 1.304322662387633e+17, 1.30432266246107e+17, 1.304322662534508e+17, 1.304322662607945e+17, 1.30432266267982e+17, 1.304322662753257e+17, 1.304322662826694e+17, 1.304322662901696e+17, 1.304322662975133e+17, 1.304322663050132e+17, 1.30432266312357e+17, 1.304322663195444e+17, 1.304322663268882e+17, 1.304322663343882e+17, 1.304322663420445e+17, 1.30432266349232e+17, 1.304322663565757e+17, 1.304322663639195e+17, 1.304322663712632e+17, 1.304322663784507e+17, 1.304322663857944e+17, 1.304322663932945e+17, 1.304322664006383e+17, 1.304322664079821e+17, 1.304322664153258e+17, 1.304322664226696e+17, 1.304322664300133e+17, 1.304322664375132e+17, 1.304322664450132e+17, 1.304322664522007e+17, 1.304322664597007e+17, 1.304322664670445e+17, 1.304322664745445e+17, 1.304322664818883e+17, 1.304322664893883e+17, 1.304322664968882e+17, 1.304322665042319e+17, 1.30432266511732e+17, 1.304322665190757e+17, 1.304322665264196e+17, 1.304322665337633e+17, 1.304322665412632e+17, 1.304322665484508e+17, 1.304322665557946e+17, 1.304322665631383e+17, 1.30432266570482e+17, 1.30432266577982e+17, 1.304322665853258e+17, 1.304322665926696e+17, 1.304322666001695e+17, 1.304322666076695e+17, 1.304322666150132e+17, 1.30432266622357e+17, 1.304322666295444e+17, 1.304322666370445e+17, 1.304322666443884e+17, 1.304322666518883e+17, 1.30432266659232e+17, 1.304322666665756e+17, 1.304322666740758e+17, 1.304322666815758e+17, 1.304322666890757e+17, 1.304322666965757e+17, 1.304322667037633e+17, 1.304322667111071e+17, 1.30432266718607e+17, 1.304322667257944e+17, 1.304322667331383e+17, 1.304322667406382e+17, 1.30432266747982e+17, 1.304322667554821e+17, 1.304322667628257e+17, 1.304322667701696e+17, 1.304322667775133e+17, 1.304322667850132e+17, 1.30432266792357e+17, 1.30432266799857e+17, 1.304322668070445e+17, 1.304322668145445e+17, 1.304322668218883e+17, 1.30432266829232e+17, 1.30432266836732e+17, 1.304322668440758e+17, 1.304322668515757e+17, 1.304322668589196e+17, 1.304322668662633e+17, 1.30432266873607e+17, 1.304322668809507e+17, 1.304322668882944e+17, 1.304322668956381e+17, 1.30432266902982e+17, 1.304322669103258e+17, 1.304322669178258e+17, 1.304322669251695e+17, 1.304322669325133e+17, 1.304322669400132e+17, 1.304322669473571e+17, 1.304322669547008e+17, 1.304322669620445e+17, 1.30432266969232e+17, 1.30432266976732e+17, 1.304322669842319e+17, 1.304322669918883e+17, 1.30432266999232e+17, 1.304322670065757e+17, 1.304322670139195e+17, 1.304322670214195e+17, 1.304322670287633e+17, 1.304322670362633e+17, 1.304322670437632e+17, 1.304322670511069e+17, 1.304322670584507e+17, 1.304322670659507e+17, 1.304322670732945e+17, 1.304322670807945e+17, 1.304322670881382e+17, 1.30432267095482e+17, 1.304322671028257e+17, 1.304322671101695e+17, 1.304322671175133e+17, 1.304322671248571e+17, 1.304322671322008e+17, 1.304322671398569e+17, 1.304322671473571e+17, 1.304322671547008e+17, 1.304322671620445e+17, 1.304322671693883e+17, 1.30432267176732e+17, 1.304322671840758e+17, 1.304322671915758e+17, 1.304322671989196e+17, 1.304322672064195e+17, 1.304322672137632e+17, 1.304322672209508e+17, 1.304322672284507e+17, 1.304322672359507e+17, 1.304322672432946e+17, 1.304322672506383e+17, 1.304322672578258e+17, 1.304322672653258e+17, 1.304322672726696e+17, 1.304322672800133e+17, 1.304322672875132e+17, 1.30432267294857e+17, 1.304322673022008e+17, 1.304322673095444e+17, 1.304322673168883e+17, 1.304322673242321e+17, 1.30432267331732e+17, 1.304322673390757e+17, 1.304322673465757e+17, 1.304322673537632e+17, 1.304322673611071e+17, 1.30432267368607e+17, 1.304322673757946e+17, 1.304322673831383e+17, 1.304322673906382e+17, 1.30432267397982e+17, 1.304322674053257e+17, 1.304322674126694e+17, 1.304322674200133e+17, 1.304322674273571e+17, 1.304322674345445e+17, 1.304322674420445e+17, 1.304322674493883e+17, 1.30432267456732e+17, 1.304322674642319e+17, 1.304322674717321e+17, 1.304322674790758e+17, 1.304322674865757e+17, 1.304322674939195e+17, 1.304322675012632e+17, 1.30432267508607e+17, 1.304322675159507e+17, 1.304322675232945e+17, 1.304322675306383e+17, 1.304322675381382e+17, 1.30432267545482e+17, 1.304322675528257e+17, 1.304322675601695e+17, 1.304322675675132e+17, 1.30432267574857e+17, 1.304322675822007e+17, 1.304322675895446e+17, 1.304322675968883e+17, 1.304322676043882e+17, 1.30432267611732e+17, 1.304322676190757e+17, 1.304322676264195e+17, 1.304322676337632e+17, 1.304322676411069e+17, 1.304322676484508e+17, 1.304322676557946e+17, 1.304322676632945e+17, 1.304322676706382e+17, 1.30432267677982e+17, 1.304322676856383e+17, 1.304322676931382e+17, 1.304322677004819e+17, 1.304322677078257e+17, 1.304322677153258e+17, 1.304322677226696e+17, 1.30432267729857e+17, 1.304322677372008e+17, 1.304322677447008e+17, 1.304322677520445e+17, 1.30432267759232e+17, 1.304322677665757e+17, 1.304322677742321e+17, 1.304322677814195e+17, 1.304322677889196e+17, 1.304322677964195e+17, 1.304322678037632e+17, 1.304322678111069e+17, 1.304322678184507e+17, 1.304322678257944e+17, 1.304322678331383e+17, 1.30432267840482e+17, 1.304322678479821e+17, 1.30432267855482e+17, 1.304322678626694e+17, 1.304322678700132e+17, 1.304322678773569e+17, 1.304322678847007e+17, 1.304322678922007e+17, 1.304322678995444e+17, 1.304322679070445e+17, 1.304322679145445e+17, 1.304322679218883e+17, 1.304322679293883e+17, 1.30432267936732e+17, 1.304322679442319e+17, 1.304322679517321e+17, 1.304322679590757e+17, 1.304322679664196e+17, 1.304322679737633e+17, 1.304322679809508e+17, 1.304322679884507e+17, 1.304322679957944e+17, 1.304322680032945e+17, 1.304322680106383e+17, 1.30432268017982e+17, 1.304322680253257e+17, 1.304322680326694e+17, 1.304322680403258e+17, 1.304322680476695e+17, 1.304322680551695e+17, 1.30432268062357e+17, 1.304322680697007e+17, 1.304322680770445e+17, 1.304322680843882e+17, 1.304322680918883e+17, 1.30432268099232e+17, 1.304322681065757e+17, 1.304322681143882e+17, 1.304322681218883e+17, 1.30432268129232e+17, 1.304322681365757e+17, 1.304322681440756e+17, 1.304322681515758e+17, 1.304322681589196e+17, 1.304322681662633e+17, 1.30432268173607e+17, 1.304322681831383e+17, 1.30432268190482e+17, 1.304322681978258e+17, 1.304322682050132e+17, 1.30432268212357e+17, 1.304322682195446e+17, 1.30432268226732e+17, 1.304322682340758e+17, 1.304322682415758e+17, 1.304322682487633e+17, 1.304322682559507e+17, 1.304322682631382e+17, 1.30432268270482e+17, 1.304322682778258e+17, 1.304322682850132e+17, 1.30432268292357e+17, 1.304322682997007e+17, 1.304322683068882e+17, 1.304322683142319e+17, 1.304322683215758e+17, 1.304322683287633e+17, 1.304322683359507e+17, 1.304322683432945e+17, 1.304322683506382e+17, 1.304322683578257e+17, 1.304322683650132e+17, 1.30432268372357e+17, 1.304322683795444e+17, 1.30432268386732e+17, 1.304322683940758e+17, 1.304322684014195e+17, 1.304322684086071e+17, 1.304322684157946e+17, 1.304322684231383e+17, 1.304322684303258e+17, 1.304322684375132e+17, 1.30432268444857e+17, 1.304322684520444e+17, 1.30432268459232e+17, 1.304322684664195e+17, 1.30432268473607e+17, 1.304322684807945e+17, 1.304322684881384e+17, 1.30432268495482e+17, 1.304322685026696e+17, 1.304322685100133e+17, 1.304322685173571e+17, 1.304322685245445e+17, 1.304322685318883e+17, 1.30432268539232e+17, 1.304322685465757e+17, 1.304322685537633e+17, 1.304322685611071e+17, 1.304322685684507e+17, 1.304322685756383e+17, 1.304322685831382e+17, 1.304322685904819e+17, 1.304322685978257e+17, 1.304322686050132e+17, 1.30432268612357e+17, 1.304322686195444e+17, 1.304322686268882e+17, 1.304322686342319e+17, 1.304322686417321e+17, 1.304322686489194e+17, 1.304322686562633e+17, 1.30432268663607e+17, 1.304322686709508e+17, 1.304322686781382e+17, 1.30432268685482e+17, 1.304322686928257e+17, 1.304322687000133e+17, 1.304322687073571e+17, 1.304322687147008e+17, 1.304322687220445e+17, 1.30432268729232e+17, 1.304322687365757e+17, 1.304322687437633e+17, 1.304322687511071e+17, 1.304322687582945e+17, 1.304322687659507e+17, 1.30432268772982e+17, 1.304322687803258e+17, 1.304322687875132e+17, 1.304322687951695e+17, 1.304322688025132e+17, 1.304322688097007e+17, 1.304322688170445e+17, 1.304322688245445e+17, 1.304322688318883e+17, 1.30432268839232e+17, 1.304322688465757e+17, 1.304322688540758e+17, 1.304322688612632e+17, 1.304322688687633e+17, 1.304322688759507e+17, 1.304322688837632e+17, 1.304322688909508e+17, 1.304322688987633e+17, 1.30432268906107e+17, 1.304322689134508e+17, 1.304322689207945e+17, 1.304322689281382e+17, 1.304322689353258e+17, 1.304322689428257e+17, 1.304322689501695e+17, 1.304322689576695e+17, 1.304322689651695e+17, 1.30432268972357e+17, 1.304322689797007e+17, 1.304322689872008e+17, 1.304322689945445e+17, 1.304322690020445e+17, 1.30432269009232e+17, 1.304322690165757e+17, 1.304322690239196e+17, 1.304322690312634e+17, 1.304322690389194e+17, 1.304322690464196e+17, 1.304322690537633e+17, 1.304322690612632e+17, 1.30432269068607e+17, 1.304322690757944e+17, 1.304322690831383e+17, 1.304322690906382e+17, 1.304322690979821e+17, 1.304322691053257e+17, 1.304322691125133e+17, 1.304322691203258e+17, 1.304322691276695e+17, 1.30432269134857e+17, 1.304322691426694e+17, 1.304322691509508e+17, 1.304322691582945e+17, 1.304322691656383e+17, 1.304322691731382e+17, 1.304322691803258e+17, 1.304322691876695e+17, 1.304322691953258e+17, 1.304322692026696e+17, 1.304322692100133e+17, 1.304322692178258e+17, 1.304322692250132e+17, 1.30432269232357e+17, 1.304322692397007e+17, 1.304322692473571e+17, 1.304322692543882e+17, 1.304322692618883e+17, 1.30432269269232e+17, 1.304322692765757e+17, 1.304322692839196e+17, 1.304322692914195e+17, 1.304322692989194e+17, 1.304322693062632e+17, 1.30432269313607e+17, 1.304322693212632e+17, 1.30432269328607e+17, 1.304322693359507e+17, 1.304322693437632e+17, 1.304322693509508e+17, 1.304322693582945e+17, 1.304322693656383e+17, 1.30432269372982e+17, 1.304322693803258e+17, 1.304322693875132e+17, 1.304322693950132e+17, 1.304322694026694e+17, 1.30432269409857e+17, 1.304322694172008e+17, 1.304322694250132e+17, 1.30432269432357e+17, 1.304322694395446e+17, 1.304322694473571e+17, 1.304322694545445e+17, 1.304322694620445e+17, 1.304322694697007e+17, 1.304322694770445e+17, 1.304322694845445e+17, 1.304322694920444e+17, 1.304322694995446e+17, 1.30432269506732e+17, 1.304322695143882e+17, 1.30432269521732e+17, 1.304322695290757e+17, 1.30432269536732e+17, 1.304322695439196e+17, 1.304322695512634e+17, 1.304322695589194e+17, 1.304322695662632e+17, 1.30432269573607e+17, 1.304322695809508e+17, 1.30432269588607e+17, 1.30432269596107e+17, 1.304322696037632e+17, 1.304322696111069e+17, 1.304322696184507e+17, 1.30432269626107e+17, 1.304322696334508e+17, 1.304322696406382e+17, 1.304322696484508e+17, 1.304322696557944e+17, 1.304322696631383e+17, 1.304322696707945e+17, 1.304322696781382e+17, 1.304322696853257e+17, 1.304322696931382e+17, 1.304322697004819e+17, 1.304322697078257e+17, 1.30432269715482e+17, 1.304322697228257e+17, 1.304322697300133e+17, 1.304322697387631e+17, 1.304322697462633e+17, 1.304322697539195e+17, 1.304322697612632e+17, 1.30432269768607e+17, 1.304322697759508e+17, 1.304322697832945e+17, 1.304322697906382e+17, 1.30432269797982e+17, 1.304322698053257e+17, 1.30432269812982e+17, 1.304322698203258e+17, 1.304322698278257e+17, 1.304322698353257e+17, 1.304322698428257e+17, 1.304322698503258e+17, 1.304322698576695e+17, 1.304322698650132e+17, 1.30432269872357e+17, 1.30432269879857e+17, 1.304322698872008e+17, 1.30432269894857e+17, 1.304322699022007e+17, 1.304322699097007e+17, 1.304322699170445e+17, 1.304322699247007e+17, 1.304322699320445e+17, 1.304322699395444e+17, 1.304322699470445e+17, 1.304322699545445e+17, 1.304322699620444e+17, 1.30432269970482e+17, 1.30432269977982e+17, 1.304322699856383e+17, 1.30432269993607e+17, 1.304322700011069e+17, 1.304322700084507e+17, 1.304322700159508e+17, 1.304322700234508e+17, 1.304322700307945e+17, 1.304322700382945e+17, 1.304322700457946e+17, 1.304322700542321e+17, 1.30432270061732e+17, 1.30432270069232e+17, 1.304322700765757e+17, 1.304322700837632e+17, 1.304322700912632e+17, 1.304322700989196e+17, 1.304322701062633e+17, 1.304322701137633e+17, 1.304322701211071e+17, 1.30432270128607e+17, 1.30432270136107e+17, 1.304322701440758e+17, 1.304322701515757e+17, 1.304322701589196e+17, 1.304322701664195e+17, 1.304322701737632e+17, 1.304322701811069e+17, 1.304322701886071e+17, 1.30432270196107e+17, 1.304322702034508e+17, 1.304322702109508e+17, 1.304322702184508e+17, 1.304322702259507e+17, 1.304322702332945e+17, 1.304322702407945e+17, 1.304322702481382e+17, 1.304322702556383e+17, 1.304322702631383e+17, 1.30432270270482e+17, 1.30432270277982e+17, 1.30432270285482e+17, 1.30432270292982e+17, 1.304322703003258e+17, 1.304322703078257e+17, 1.304322703153257e+17, 1.304322703228257e+17, 1.304322703301696e+17, 1.304322703376695e+17, 1.304322703453258e+17, 1.304322703532945e+17, 1.304322703607944e+17, 1.304322703681382e+17, 1.304322703756383e+17, 1.304322703831383e+17, 1.304322703907945e+17, 1.304322703981382e+17, 1.304322704056383e+17, 1.304322704132945e+17, 1.304322704206382e+17, 1.304322704284508e+17, 1.304322704359507e+17, 1.30432270443607e+17, 1.304322704511069e+17, 1.304322704589196e+17, 1.304322704662633e+17, 1.30432270473607e+17, 1.304322704812632e+17, 1.304322704884507e+17, 1.304322704959508e+17, 1.304322705034508e+17, 1.304322705109508e+17, 1.304322705181382e+17, 1.304322705257946e+17, 1.304322705331383e+17, 1.30432270540482e+17, 1.304322705482945e+17, 1.30432270555482e+17, 1.304322705628257e+17, 1.304322705704819e+17, 1.304322705778258e+17, 1.304322705851695e+17, 1.30432270592982e+17, 1.304322706003258e+17, 1.304322706076695e+17, 1.304322706153257e+17, 1.304322706226694e+17, 1.304322706300132e+17, 1.304322706376695e+17, 1.304322706450132e+17, 1.30432270652357e+17, 1.30432270659857e+17, 1.304322706672008e+17, 1.304322706745445e+17, 1.304322706822007e+17, 1.304322706897007e+17, 1.304322706970445e+17, 1.304322707045445e+17, 1.304322707120445e+17, 1.304322707193883e+17, 1.304322707268882e+17, 1.304322707343882e+17, 1.30432270741732e+17, 1.304322707493883e+17, 1.304322707568882e+17, 1.304322707645445e+17, 1.304322707718883e+17, 1.30432270779232e+17, 1.304322707868883e+17, 1.304322707943882e+17, 1.30432270801732e+17, 1.304322708093883e+17, 1.304322708165757e+17, 1.304322708239195e+17, 1.304322708312632e+17, 1.30432270838607e+17, 1.304322708459507e+17, 1.304322708532945e+17, 1.30432270860482e+17, 1.304322708678258e+17, 1.304322708751695e+17, 1.304322708825133e+17, 1.304322708900132e+17, 1.304322708975133e+17, 1.304322709048571e+17, 1.304322709120445e+17, 1.304322709193883e+17, 1.30432270926732e+17, 1.304322709340758e+17, 1.304322709415757e+17, 1.304322709489194e+17, 1.304322709564196e+17, 1.304322709639195e+17, 1.304322709709508e+17, 1.304322709782945e+17, 1.304322709856383e+17, 1.30432270992982e+17, 1.304322710004819e+17, 1.304322710078257e+17, 1.30432271015482e+17, 1.304322710228257e+17, 1.304322710301695e+17, 1.304322710378258e+17, 1.304322710451695e+17, 1.304322710665757e+17, 1.304322710743882e+17, 1.30432271081732e+17, 1.304322710890757e+17, 1.304322710965757e+17, 1.304322711039195e+17, 1.304322711112634e+17, 1.304322711190757e+17, 1.304322711264196e+17, 1.304322711337633e+17, 1.304322711414195e+17, 1.304322711487631e+17, 1.304322711562633e+17, 1.304322711637633e+17, 1.304322711711071e+17, 1.304322711784507e+17, 1.30432271186107e+17, 1.30432271193607e+17, 1.304322712009508e+17, 1.304322712084508e+17, 1.304322712159507e+17, 1.304322712232945e+17, 1.304322712307945e+17, 1.304322712395444e+17, 1.304322712472008e+17, 1.304322712550132e+17, 1.304322712628257e+17, 1.304322712714195e+17, 1.304322712787633e+17, 1.304322712862633e+17, 1.304322712937632e+17, 1.304322713012632e+17, 1.30432271308607e+17, 1.30432271316107e+17, 1.304322713234508e+17, 1.304322713306383e+17, 1.304322713379821e+17, 1.304322713453258e+17, 1.304322713526696e+17, 1.304322713606382e+17, 1.304322713681382e+17, 1.304322713756383e+17, 1.304322713831383e+17, 1.30432271390482e+17, 1.304322713979821e+17, 1.304322714053258e+17, 1.304322714126696e+17, 1.304322714200133e+17, 1.304322714273571e+17, 1.304322714345445e+17, 1.304322714422007e+17, 1.304322714495444e+17, 1.304322714567319e+17, 1.304322714642321e+17, 1.304322714715758e+17, 1.30432271479232e+17, 1.30432271486732e+17, 1.304322714942321e+17, 1.304322715015757e+17, 1.304322715089196e+17, 1.304322715162633e+17, 1.304322715234508e+17, 1.304322715307945e+17, 1.304322715381382e+17, 1.304322715456383e+17, 1.30432271552982e+17, 1.304322715603258e+17, 1.304322715678257e+17, 1.304322715751694e+17, 1.304322715825132e+17, 1.304322715903256e+17, 1.304322715978258e+17, 1.304322716051695e+17, 1.304322716125133e+17, 1.30432271619857e+17, 1.304322716273571e+17, 1.304322716350132e+17, 1.30432271642357e+17, 1.30432271649857e+17, 1.304322716572008e+17, 1.304322716647008e+17, 1.304322716722007e+17, 1.304322716793883e+17, 1.304322716868882e+17, 1.304322716942319e+17, 1.304322717022007e+17, 1.304322717093882e+17, 1.30432271719232e+17, 1.304322717275132e+17, 1.304322717347008e+17, 1.304322717428257e+17, 1.304322717501695e+17, 1.304322717575132e+17, 1.30432271764857e+17, 1.304322717722008e+17, 1.304322717795446e+17, 1.304322717873571e+17, 1.304322717947008e+17, 1.304322718020445e+17, 1.304322718095444e+17, 1.304322718170445e+17, 1.304322718240758e+17, 1.304322718314195e+17, 1.30432271839232e+17, 1.304322718462633e+17, 1.30432271853607e+17, 1.304322718609508e+17, 1.30432271868607e+17, 1.304322718757944e+17, 1.304322718831382e+17, 1.304322718907945e+17, 1.304322718982944e+17, 1.30432271905482e+17, 1.304322719132945e+17, 1.304322719206383e+17, 1.304322719278258e+17, 1.30432271935482e+17, 1.30432271942982e+17, 1.304322719503258e+17, 1.304322719587633e+17, 1.30432271966107e+17, 1.304322719734508e+17, 1.304322719811069e+17, 1.304322719884508e+17, 1.304322719959507e+17, 1.304322720032945e+17, 1.304322720107945e+17, 1.30432272017982e+17, 1.304322720253257e+17, 1.304322720331382e+17, 1.304322720403258e+17, 1.304322720478257e+17, 1.30432272055482e+17, 1.304322720628257e+17, 1.304322720701695e+17, 1.304322720778258e+17, 1.304322720851695e+17, 1.30432272092357e+17, 1.304322721001695e+17, 1.304322721075132e+17, 1.304322721148571e+17, 1.304322721225133e+17, 1.30432272129857e+17, 1.304322721372008e+17, 1.30432272144857e+17, 1.30432272152357e+17, 1.304322721601695e+17, 1.304322721675132e+17, 1.304322721751695e+17, 1.304322721825133e+17, 1.30432272189857e+17, 1.304322721989196e+17, 1.30432272206732e+17, 1.304322722139196e+17, 1.304322722218883e+17, 1.30432272229232e+17, 1.304322722364196e+17, 1.30432272243607e+17, 1.304322722511071e+17, 1.304322722582945e+17, 1.304322722657944e+17, 1.30432272272982e+17, 1.304322722803258e+17, 1.304322722876695e+17, 1.304322722950132e+17, 1.30432272302357e+17, 1.304322723097007e+17, 1.304322723175132e+17, 1.30432272324857e+17, 1.304322723322007e+17, 1.30432272339857e+17, 1.304322723472008e+17, 1.304322723545445e+17, 1.304322723620445e+17, 1.304322723693883e+17, 1.304322723765757e+17, 1.304322723839195e+17, 1.304322723912632e+17, 1.30432272398607e+17, 1.304322724059507e+17, 1.304322724132945e+17, 1.30432272420482e+17, 1.304322724278258e+17, 1.30432272435482e+17, 1.304322724434508e+17, 1.304322724507945e+17, 1.304322724582945e+17, 1.304322724656383e+17, 1.30432272472982e+17, 1.304322724803256e+17, 1.304322724879821e+17, 1.304322724953258e+17, 1.304322725028257e+17, 1.30432272510482e+17, 1.304322725176695e+17, 1.304322725250132e+17, 1.30432272532357e+17, 1.30432272539857e+17, 1.304322725472008e+17, 1.304322725551695e+17, 1.304322725626696e+17, 1.304322725700133e+17, 1.304322725773571e+17, 1.304322725847008e+17, 1.304322725920444e+17, 1.30432272599857e+17, 1.304322726072008e+17, 1.304322726145445e+17, 1.304322726220445e+17, 1.304322726293883e+17, 1.304322726365757e+17, 1.304322726439195e+17, 1.304322726512632e+17, 1.30432272658607e+17, 1.304322726659507e+17, 1.304322726743884e+17, 1.30432272682982e+17, 1.304322726903258e+17, 1.304322726984507e+17, 1.304322727056383e+17, 1.304322727131382e+17, 1.30432272720482e+17, 1.304322727276695e+17, 1.304322727351695e+17, 1.304322727425133e+17, 1.304322727501695e+17, 1.304322727573569e+17, 1.304322727647007e+17, 1.304322727725133e+17, 1.30432272779857e+17, 1.304322727870445e+17, 1.304322727950132e+17, 1.30432272802982e+17, 1.304322728103258e+17, 1.304322728175132e+17, 1.304322728251695e+17, 1.304322728325133e+17, 1.304322728401695e+17, 1.304322728476695e+17, 1.304322728550132e+17, 1.304322728626696e+17, 1.304322728700133e+17, 1.304322728775132e+17, 1.30432272884857e+17, 1.30432272892357e+17, 1.30432272899857e+17, 1.304322729070446e+17, 1.304322729150132e+17, 1.304322729222008e+17, 1.304322729295446e+17, 1.304322729370445e+17, 1.304322729443882e+17, 1.304322729518883e+17, 1.30432272959232e+17, 1.304322729665757e+17, 1.304322729739195e+17, 1.304322729812632e+17, 1.304322729884508e+17, 1.304322729957946e+17, 1.304322730032945e+17, 1.30432273010482e+17, 1.304322730182945e+17, 1.304322730256383e+17, 1.30432273032982e+17, 1.304322730406382e+17, 1.304322730481382e+17, 1.30432273055482e+17, 1.304322730628257e+17, 1.304322730701695e+17, 1.304322730775132e+17, 1.304322730851695e+17, 1.304322730926694e+17, 1.304322731000132e+17, 1.304322731075133e+17, 1.304322731148571e+17, 1.304322731222008e+17, 1.304322731300133e+17, 1.304322731372008e+17, 1.304322731445445e+17, 1.304322731532945e+17, 1.304322731609508e+17, 1.30432273168607e+17, 1.304322731759507e+17, 1.304322731832945e+17, 1.304322731907945e+17, 1.304322731981382e+17, 1.30432273205482e+17, 1.304322732132946e+17, 1.30432273220482e+17, 1.304322732278258e+17, 1.30432273235482e+17, 1.30432273242982e+17, 1.304322732503258e+17, 1.30432273257982e+17, 1.304322732653257e+17, 1.304322732728257e+17, 1.30432273280482e+17, 1.304322732876695e+17, 1.304322732950132e+17, 1.304322733025133e+17, 1.30432273309857e+17, 1.304322733170445e+17, 1.30432273324857e+17, 1.304322733322007e+17, 1.304322733395446e+17, 1.304322733472008e+17, 1.304322733547008e+17, 1.304322733620445e+17, 1.304322733695444e+17, 1.304322733768883e+17, 1.304322733842321e+17, 1.304322733925133e+17, 1.304322734001695e+17, 1.304322734073571e+17, 1.30432273414857e+17, 1.304322734222008e+17, 1.304322734295444e+17, 1.304322734368883e+17, 1.304322734447008e+17, 1.304322734522007e+17, 1.304322734595444e+17, 1.304322734670445e+17, 1.304322734745445e+17, 1.304322734818883e+17, 1.304322734893882e+17, 1.304322734967319e+17, 1.304322735042321e+17, 1.304322735120445e+17, 1.304322735195446e+17, 1.30432273526732e+17, 1.304322735342321e+17, 1.304322735415757e+17, 1.304322735489196e+17, 1.304322735564195e+17, 1.304322735637633e+17, 1.304322735711071e+17, 1.304322735784508e+17, 1.304322735856383e+17, 1.30432273592982e+17, 1.304322736003258e+17, 1.304322736076695e+17, 1.304322736150132e+17, 1.30432273622357e+17, 1.304322736332945e+17, 1.304322736418883e+17, 1.30432273649232e+17, 1.304322736575132e+17, 1.30432273664857e+17, 1.304322736722007e+17, 1.304322736795444e+17, 1.30432273686732e+17, 1.304322736940756e+17, 1.304322737015757e+17, 1.304322737089196e+17, 1.304322737161069e+17, 1.304322737234508e+17, 1.304322737312632e+17, 1.304322737384508e+17, 1.304322737457944e+17, 1.304322737534508e+17, 1.304322737607945e+17, 1.304322737681382e+17, 1.304322737759507e+17, 1.304322737832945e+17, 1.30432273790482e+17, 1.304322737982945e+17, 1.304322738057944e+17, 1.304322738137632e+17, 1.304322738209508e+17, 1.304322738287633e+17, 1.30432273836107e+17, 1.304322738434508e+17, 1.304322738509507e+17, 1.304322738582945e+17, 1.304322738656383e+17, 1.304322738739195e+17, 1.304322738815758e+17, 1.304322738889196e+17, 1.304322738968883e+17, 1.304322739039195e+17, 1.304322739112632e+17, 1.30432273918607e+17, 1.304322739262633e+17, 1.304322739336069e+17, 1.304322739407945e+17, 1.30432273948607e+17, 1.304322739559507e+17, 1.304322739632945e+17, 1.304322739709508e+17, 1.304322739781384e+17, 1.304322739854821e+17, 1.304322739932946e+17, 1.304322740009507e+17, 1.304322740082944e+17, 1.304322740157946e+17, 1.30432274022982e+17, 1.304322740303258e+17, 1.304322740378258e+17, 1.304322740451695e+17, 1.304322740526694e+17, 1.304322740601695e+17, 1.304322740675132e+17, 1.30432274074857e+17, 1.304322740822007e+17, 1.304322740895444e+17, 1.304322740968882e+17, 1.304322741042319e+17, 1.304322741126694e+17, 1.304322741201695e+17, 1.304322741273569e+17, 1.304322741353257e+17, 1.304322741426696e+17, 1.304322741500133e+17, 1.304322741579821e+17, 1.304322741653258e+17, 1.304322741726696e+17, 1.304322741800133e+17, 1.304322741872008e+17, 1.304322741947008e+17, 1.304322742025133e+17, 1.30432274209857e+17, 1.304322742172008e+17, 1.304322742247008e+17, 1.30432274232357e+17, 1.304322742397007e+17, 1.304322742470445e+17, 1.304322742543882e+17, 1.304322742618883e+17, 1.304322742695444e+17, 1.304322742768882e+17, 1.304322742840756e+17, 1.304322742914194e+17, 1.304322742990757e+17, 1.304322743062633e+17, 1.30432274313607e+17, 1.30432274321732e+17, 1.304322743290757e+17, 1.304322743364195e+17, 1.304322743437633e+17, 1.304322743514195e+17, 1.304322743587633e+17, 1.30432274366107e+17, 1.30432274373607e+17, 1.304322743812632e+17, 1.30432274388607e+17, 1.304322743959507e+17, 1.30432274403607e+17, 1.304322744109508e+17, 1.304322744182944e+17, 1.304322744259508e+17, 1.304322744331383e+17, 1.30432274440482e+17, 1.304322744482945e+17, 1.304322744556383e+17, 1.30432274462982e+17, 1.30432274470482e+17, 1.30432274477982e+17, 1.304322744851695e+17, 1.30432274492982e+17, 1.304322745003258e+17, 1.304322745076695e+17, 1.304322745151695e+17, 1.304322745225133e+17, 1.30432274529857e+17, 1.304322745372008e+17, 1.304322745448571e+17, 1.30432274552357e+17, 1.304322745600133e+17, 1.304322745672006e+17, 1.304322745745445e+17, 1.304322745822008e+17, 1.304322745912632e+17, 1.304322745989196e+17, 1.304322746067319e+17, 1.304322746143882e+17, 1.30432274621732e+17, 1.304322746290757e+17, 1.304322746364195e+17, 1.304322746437632e+17, 1.304322746514195e+17, 1.304322746587633e+17, 1.304322746662632e+17, 1.304322746737633e+17, 1.304322746811071e+17, 1.30432274688607e+17, 1.30432274696107e+17, 1.30432274703607e+17, 1.304322747115757e+17, 1.304322747189194e+17, 1.304322747264195e+17, 1.304322747339196e+17, 1.304322747414195e+17, 1.304322747489194e+17, 1.304322747562633e+17, 1.30432274763607e+17, 1.304322747711071e+17, 1.304322747784508e+17, 1.304322747857944e+17, 1.304322747934508e+17, 1.304322748009508e+17, 1.304322748082945e+17, 1.304322748159507e+17, 1.304322748232945e+17, 1.304322748312632e+17, 1.30432274838607e+17, 1.304322748459507e+17, 1.30432274853607e+17, 1.304322748607945e+17, 1.304322748681384e+17, 1.304322748754821e+17, 1.304322748828257e+17, 1.304322748901695e+17, 1.304322748975132e+17, 1.304322749051695e+17, 1.304322749125133e+17, 1.30432274919857e+17, 1.304322749272008e+17, 1.304322749345445e+17, 1.304322749420444e+17, 1.304322749500132e+17, 1.304322749573571e+17, 1.304322749647008e+17, 1.30432274972357e+17, 1.30432274979857e+17, 1.304322749872008e+17, 1.30432274994857e+17, 1.304322750028257e+17, 1.304322750103258e+17, 1.30432275017982e+17, 1.304322750254821e+17, 1.304322750332946e+17, 1.304322750406383e+17, 1.304322750481382e+17, 1.304322750556381e+17, 1.30432275062982e+17, 1.304322750718883e+17, 1.304322750793882e+17, 1.30432275086732e+17, 1.304322750945444e+17, 1.30432275102357e+17, 1.30432275109857e+17, 1.304322751172008e+17, 1.30432275124857e+17, 1.304322751326696e+17, 1.304322751401695e+17, 1.304322751476695e+17, 1.304322751551695e+17, 1.304322751626696e+17, 1.304322751701695e+17, 1.304322751775132e+17, 1.304322751850132e+17, 1.304322751925133e+17, 1.304322752000132e+17, 1.30432275207982e+17, 1.30432275215482e+17, 1.30432275222982e+17, 1.304322752304819e+17, 1.304322752376695e+17, 1.304322752450132e+17, 1.304322752525132e+17, 1.304322752601695e+17, 1.304322752675132e+17, 1.30432275274857e+17, 1.30432275282357e+17, 1.30432275289857e+17, 1.304322752973571e+17, 1.304322753048571e+17, 1.304322753131383e+17, 1.304322753211069e+17, 1.30432275328607e+17, 1.30432275336107e+17, 1.304322753434508e+17, 1.304322753507945e+17, 1.304322753581382e+17, 1.30432275365482e+17, 1.304322753728257e+17, 1.304322753801695e+17, 1.304322753878257e+17, 1.304322753948571e+17, 1.304322754022008e+17, 1.304322754095444e+17, 1.304322754172008e+17, 1.304322754245445e+17, 1.304322754322007e+17, 1.304322754395444e+17, 1.304322754468882e+17, 1.304322754543882e+17, 1.304322754618883e+17, 1.304322754690757e+17, 1.304322754764195e+17, 1.304322754840758e+17, 1.30432275491732e+17, 1.304322754990757e+17, 1.304322755065757e+17, 1.304322755139196e+17, 1.304322755211071e+17, 1.304322755289194e+17, 1.304322755362633e+17, 1.304322755434508e+17, 1.304322755532945e+17, 1.304322755620444e+17, 1.304322755695444e+17, 1.304322755782945e+17, 1.304322755857944e+17, 1.304322755932945e+17, 1.304322756006382e+17, 1.304322756079821e+17, 1.304322756153258e+17, 1.304322756226696e+17, 1.30432275630482e+17, 1.304322756378258e+17, 1.304322756451695e+17, 1.304322756528257e+17, 1.304322756601695e+17, 1.304322756675132e+17, 1.304322756753257e+17, 1.304322756826694e+17, 1.304322756900133e+17, 1.304322756973571e+17, 1.30432275704857e+17, 1.30432275712357e+17, 1.304322757197007e+17, 1.304322757268882e+17, 1.304322757342319e+17, 1.304322757415757e+17, 1.304322757489196e+17, 1.304322757564196e+17, 1.304322757639195e+17, 1.304322757711071e+17, 1.30432275778607e+17, 1.304322757859507e+17, 1.304322757937632e+17, 1.304322758012632e+17, 1.304322758087633e+17, 1.304322758164196e+17, 1.30432275823607e+17, 1.304322758307945e+17, 1.304322758381382e+17, 1.304322758456383e+17, 1.304322758531382e+17, 1.304322758603258e+17, 1.304322758681382e+17, 1.304322758753258e+17, 1.304322758826696e+17, 1.304322758900133e+17, 1.30432275898607e+17, 1.304322759057946e+17, 1.30432275913607e+17, 1.304322759211071e+17, 1.304322759284508e+17, 1.304322759357944e+17, 1.304322759431383e+17, 1.304322759504819e+17, 1.304322759578257e+17, 1.304322759651695e+17, 1.304322759725133e+17, 1.30432275979857e+17, 1.304322759872008e+17, 1.304322759945445e+17, 1.304322760023571e+17, 1.304322760097007e+17, 1.304322760168883e+17, 1.304322760245444e+17, 1.30432276032982e+17, 1.304322760407945e+17, 1.304322760481382e+17, 1.30432276056107e+17, 1.304322760634508e+17, 1.304322760711071e+17, 1.304322760784508e+17, 1.304322760857944e+17, 1.304322760931383e+17, 1.304322761007945e+17, 1.304322761079821e+17, 1.304322761153257e+17, 1.304322761226696e+17, 1.304322761300133e+17, 1.304322761373571e+17, 1.304322761445445e+17, 1.304322761525133e+17, 1.30432276159857e+17, 1.304322761672008e+17, 1.304322761750132e+17, 1.304322761822008e+17, 1.304322761895446e+17, 1.304322761970445e+17, 1.304322762045445e+17, 1.304322762120445e+17, 1.304322762195444e+17, 1.304322762268882e+17, 1.304322762342319e+17, 1.304322762420444e+17, 1.304322762493883e+17, 1.30432276256732e+17, 1.304322762640758e+17, 1.30432276272357e+17, 1.304322762797007e+17, 1.304322762870445e+17, 1.30432276294857e+17, 1.304322763028257e+17, 1.304322763100132e+17, 1.304322763173569e+17, 1.304322763247007e+17, 1.30432276332357e+17, 1.304322763393883e+17, 1.30432276346732e+17, 1.304322763540758e+17, 1.304322763615758e+17, 1.304322763687633e+17, 1.30432276376107e+17, 1.304322763834508e+17, 1.304322763909508e+17, 1.30432276398607e+17, 1.304322764064195e+17, 1.30432276413607e+17, 1.304322764209508e+17, 1.30432276428607e+17, 1.304322764359507e+17, 1.304322764434508e+17, 1.304322764509508e+17, 1.304322764584507e+17, 1.304322764657946e+17, 1.304322764732945e+17, 1.304322764807945e+17, 1.304322764881382e+17, 1.304322764959507e+17, 1.304322765034508e+17, 1.30432276512982e+17, 1.304322765209507e+17, 1.304322765282945e+17, 1.304322765367319e+17, 1.304322765445444e+17, 1.304322765526696e+17, 1.304322765601695e+17, 1.304322765676695e+17, 1.304322765750132e+17, 1.30432276582982e+17, 1.304322765903258e+17, 1.304322765978258e+17, 1.30432276605482e+17, 1.30432276612982e+17, 1.304322766203258e+17, 1.304322766276695e+17, 1.30432276635482e+17, 1.304322766440758e+17, 1.304322766515757e+17, 1.304322766589194e+17, 1.304322766662633e+17, 1.30432276673607e+17, 1.304322766809508e+17, 1.304322766882945e+17, 1.304322766957944e+17, 1.304322767031382e+17, 1.304322767104819e+17, 1.304322767178257e+17, 1.304322767251695e+17, 1.304322767325133e+17, 1.304322767397007e+17, 1.304322767470445e+17, 1.304322767551695e+17, 1.304322767628257e+17, 1.304322767701696e+17, 1.304322767781382e+17, 1.30432276785482e+17, 1.304322767926696e+17, 1.304322768000133e+17, 1.304322768076695e+17, 1.304322768147008e+17, 1.304322768222007e+17, 1.304322768295444e+17, 1.304322768368882e+17, 1.304322768442321e+17, 1.304322768515758e+17, 1.304322768593883e+17, 1.304322768665757e+17, 1.304322768743882e+17, 1.30432276881732e+17, 1.304322768890757e+17, 1.304322768965757e+17, 1.304322769039195e+17, 1.304322769114195e+17, 1.304322769187633e+17, 1.304322769264195e+17, 1.304322769337632e+17, 1.304322769411069e+17, 1.30432276948607e+17, 1.304322769559507e+17, 1.304322769634508e+17, 1.304322769709508e+17, 1.304322769782944e+17, 1.30432276985482e+17, 1.304322769940756e+17, 1.304322770017321e+17, 1.304322770090757e+17, 1.304322770168883e+17, 1.304322770240758e+17, 1.304322770314195e+17, 1.30432277038607e+17, 1.30432277046107e+17, 1.304322770534508e+17, 1.304322770607945e+17, 1.304322770681382e+17, 1.30432277075482e+17, 1.304322770828257e+17, 1.304322770901695e+17, 1.304322770973569e+17, 1.304322771051695e+17, 1.304322771126694e+17, 1.304322771201696e+17, 1.304322771276695e+17, 1.304322771348571e+17, 1.30432277142357e+17, 1.304322771497007e+17, 1.304322771572008e+17, 1.304322771645445e+17, 1.30432277172357e+17, 1.304322771797007e+17, 1.304322771870445e+17, 1.304322771943882e+17, 1.304322772018883e+17, 1.304322772093883e+17, 1.30432277216732e+17, 1.304322772240758e+17, 1.304322772322007e+17, 1.30432277239857e+17, 1.304322772472008e+17, 1.30432277254857e+17, 1.30432277262357e+17, 1.304322772697007e+17, 1.304322772770445e+17, 1.304322772843882e+17, 1.30432277291732e+17, 1.304322772993883e+17, 1.30432277306732e+17, 1.304322773143882e+17, 1.30432277321732e+17, 1.304322773289194e+17, 1.30432277336732e+17, 1.304322773440758e+17, 1.304322773515758e+17, 1.304322773589196e+17, 1.304322773662633e+17, 1.30432277373607e+17, 1.304322773812632e+17, 1.304322773886071e+17, 1.304322773959508e+17, 1.304322774037633e+17, 1.304322774112632e+17, 1.304322774184508e+17, 1.304322774259507e+17, 1.304322774332945e+17, 1.304322774406382e+17, 1.304322774482945e+17, 1.304322774557944e+17, 1.304322774631382e+17, 1.304322774737633e+17, 1.304322774818883e+17, 1.30432277489232e+17, 1.304322774978257e+17, 1.304322775053258e+17, 1.304322775128257e+17, 1.304322775200133e+17, 1.304322775275132e+17, 1.304322775350132e+17, 1.304322775422007e+17, 1.304322775493883e+17, 1.304322775568883e+17, 1.304322775642321e+17, 1.304322775715758e+17, 1.304322775789196e+17, 1.304322775864195e+17, 1.304322775940758e+17, 1.304322776014195e+17, 1.304322776087633e+17, 1.304322776162632e+17, 1.304322776236069e+17, 1.304322776311071e+17, 1.304322776384508e+17, 1.304322776456383e+17, 1.304322776534508e+17, 1.304322776609508e+17, 1.304322776681382e+17, 1.304322776757944e+17, 1.304322776831382e+17, 1.30432277690482e+17, 1.304322776981382e+17, 1.30432277705482e+17, 1.30432277713607e+17, 1.304322777212632e+17, 1.30432277728607e+17, 1.304322777362633e+17, 1.30432277743607e+17, 1.304322777509508e+17, 1.304322777582944e+17, 1.304322777656383e+17, 1.304322777732945e+17, 1.304322777806383e+17, 1.304322777879821e+17, 1.304322777956383e+17, 1.30432277802982e+17, 1.30432277810482e+17, 1.304322778178258e+17, 1.304322778253257e+17, 1.304322778326696e+17, 1.304322778404819e+17, 1.304322778479821e+17, 1.304322778557946e+17, 1.30432277862982e+17, 1.304322778703258e+17, 1.304322778776695e+17, 1.30432277884857e+17, 1.30432277892357e+17, 1.304322778997007e+17, 1.304322779073571e+17, 1.304322779147008e+17, 1.304322779222008e+17, 1.30432277929857e+17, 1.304322779372008e+17, 1.304322779445445e+17, 1.304322779528257e+17, 1.304322779606382e+17, 1.304322779678258e+17, 1.304322779751695e+17, 1.304322779826694e+17, 1.30432277989857e+17, 1.304322779972008e+17, 1.304322780050132e+17, 1.304322780125133e+17, 1.30432278019857e+17, 1.304322780272008e+17, 1.304322780345445e+17, 1.304322780422007e+17, 1.304322780497007e+17, 1.304322780570445e+17, 1.304322780643882e+17, 1.304322780725132e+17, 1.304322780800133e+17, 1.304322780875132e+17, 1.30432278094857e+17, 1.304322781025133e+17, 1.30432278109857e+17, 1.304322781172008e+17, 1.304322781247008e+17, 1.304322781320444e+17, 1.304322781393882e+17, 1.304322781470445e+17, 1.304322781545445e+17, 1.304322781620445e+17, 1.304322781693883e+17, 1.304322781765757e+17, 1.304322781839196e+17, 1.304322781917321e+17, 1.304322781990758e+17, 1.304322782065757e+17, 1.304322782145445e+17, 1.30432278222357e+17, 1.304322782295446e+17, 1.304322782368883e+17, 1.304322782447008e+17, 1.304322782520445e+17, 1.304322782595444e+17, 1.304322782668882e+17, 1.304322782742319e+17, 1.304322782815757e+17, 1.304322782893883e+17, 1.304322782965757e+17, 1.304322783039195e+17, 1.30432278311732e+17, 1.304322783189196e+17, 1.304322783262633e+17, 1.304322783339196e+17, 1.304322783412634e+17, 1.304322783487633e+17, 1.304322783564196e+17, 1.30432278363607e+17, 1.304322783709508e+17, 1.304322783782945e+17, 1.304322783857944e+17, 1.30432278392982e+17, 1.304322784003258e+17, 1.304322784076695e+17, 1.304322784151695e+17, 1.304322784225133e+17, 1.304322784322007e+17, 1.304322784400132e+17, 1.304322784473569e+17, 1.304322784551695e+17, 1.304322784625133e+17, 1.304322784700133e+17, 1.304322784773571e+17, 1.304322784847008e+17, 1.304322784925133e+17, 1.30432278499857e+17, 1.304322785072008e+17, 1.304322785147007e+17, 1.30432278522357e+17, 1.304322785295446e+17, 1.304322785370445e+17, 1.304322785443882e+17, 1.304322785520445e+17, 1.304322785595444e+17, 1.304322785668883e+17, 1.304322785740758e+17, 1.304322785812632e+17, 1.304322785887633e+17, 1.304322785959507e+17, 1.304322786034508e+17, 1.304322786107945e+17, 1.304322786182945e+17, 1.304322786256383e+17, 1.304322786328259e+17, 1.304322786401696e+17, 1.304322786475133e+17, 1.304322786548571e+17, 1.304322786625133e+17, 1.30432278670482e+17, 1.304322786778258e+17, 1.304322786853257e+17, 1.304322786926694e+17, 1.304322787000132e+17, 1.304322787078258e+17, 1.304322787151695e+17, 1.304322787225133e+17, 1.304322787301695e+17, 1.304322787373571e+17, 1.304322787447008e+17, 1.304322787525133e+17, 1.30432278759857e+17, 1.304322787672008e+17, 1.304322787747007e+17, 1.304322787822008e+17, 1.30432278789857e+17, 1.304322787973571e+17, 1.304322788051694e+17, 1.304322788126696e+17, 1.304322788200133e+17, 1.304322788275132e+17, 1.30432278834857e+17, 1.304322788422007e+17, 1.304322788500133e+17, 1.304322788575132e+17, 1.304322788650132e+17, 1.30432278872357e+17, 1.304322788797007e+17, 1.304322788870445e+17, 1.304322788947008e+17, 1.304322789020445e+17, 1.304322789109508e+17, 1.304322789184508e+17, 1.304322789257944e+17, 1.304322789334508e+17, 1.304322789406382e+17, 1.30432278947982e+17, 1.304322789554821e+17, 1.30432278962982e+17, 1.304322789703256e+17, 1.304322789778258e+17, 1.304322789851695e+17, 1.304322789925133e+17, 1.304322790001695e+17, 1.304322790076695e+17, 1.304322790150132e+17, 1.304322790226694e+17, 1.304322790300132e+17, 1.304322790373571e+17, 1.30432279044857e+17, 1.304322790522007e+17, 1.304322790597007e+17, 1.304322790673571e+17, 1.304322790747008e+17, 1.304322790820444e+17, 1.304322790895444e+17, 1.304322790968883e+17, 1.304322791042321e+17, 1.304322791115758e+17, 1.304322791189196e+17, 1.304322791262633e+17, 1.304322791334508e+17, 1.304322791409508e+17, 1.30432279149232e+17, 1.304322791568882e+17, 1.304322791642319e+17, 1.304322791715757e+17, 1.304322791789196e+17, 1.304322791862633e+17, 1.30432279193607e+17, 1.304322792014195e+17, 1.304322792087633e+17, 1.30432279216107e+17, 1.304322792234508e+17, 1.304322792307945e+17, 1.304322792379821e+17, 1.304322792453258e+17, 1.304322792528257e+17, 1.304322792601695e+17, 1.304322792682945e+17, 1.304322792759507e+17, 1.304322792832945e+17, 1.30432279290482e+17, 1.304322792979821e+17, 1.304322793051695e+17, 1.304322793125133e+17, 1.30432279319857e+17, 1.304322793272008e+17, 1.304322793345445e+17, 1.304322793420444e+17, 1.304322793495444e+17, 1.304322793570445e+17, 1.304322793643884e+17, 1.304322793720445e+17, 1.304322793793883e+17, 1.304322793890757e+17, 1.30432279396732e+17, 1.304322794045445e+17, 1.30432279412982e+17, 1.304322794207945e+17, 1.304322794281382e+17, 1.30432279435482e+17, 1.304322794431383e+17, 1.304322794506383e+17, 1.304322794584508e+17, 1.30432279465482e+17, 1.304322794728257e+17, 1.304322794801695e+17, 1.304322794876695e+17, 1.304322794950132e+17, 1.30432279502357e+17, 1.304322795101695e+17, 1.304322795173571e+17, 1.304322795247008e+17, 1.304322795325133e+17, 1.30432279539857e+17, 1.304322795472008e+17, 1.304322795547007e+17, 1.304322795623571e+17, 1.304322795695446e+17, 1.304322795770445e+17, 1.304322795845444e+17, 1.304322795918883e+17, 1.304322795995444e+17, 1.304322796068883e+17, 1.304322796142321e+17, 1.304322796218883e+17, 1.304322796293883e+17, 1.304322796372008e+17, 1.304322796442321e+17, 1.304322796515758e+17, 1.304322796590757e+17, 1.304322796665757e+17, 1.304322796737632e+17, 1.304322796809508e+17, 1.304322796882944e+17, 1.304322796956383e+17, 1.30432279702982e+17, 1.30432279710482e+17, 1.304322797176695e+17, 1.30432279725482e+17, 1.304322797328257e+17, 1.304322797400133e+17, 1.304322797478258e+17, 1.304322797553257e+17, 1.304322797626694e+17, 1.304322797700133e+17, 1.304322797773571e+17, 1.304322797847008e+17, 1.304322797925133e+17, 1.304322797997007e+17, 1.304322798072008e+17, 1.304322798147007e+17, 1.304322798222007e+17, 1.304322798295446e+17, 1.304322798370445e+17, 1.304322798443882e+17, 1.30432279851732e+17, 1.304322798595444e+17, 1.304322798676695e+17, 1.304322798756383e+17, 1.304322798831383e+17, 1.304322798907945e+17, 1.304322798981382e+17, 1.30432279905482e+17, 1.304322799128257e+17, 1.304322799203258e+17, 1.304322799276695e+17, 1.304322799350132e+17, 1.304322799428257e+17, 1.304322799501695e+17, 1.304322799576695e+17, 1.304322799650132e+17, 1.304322799723571e+17, 1.304322799797009e+17, 1.304322799876695e+17, 1.304322799954821e+17, 1.304322800028257e+17, 1.304322800104819e+17, 1.304322800178258e+17, 1.304322800250132e+17, 1.30432280032357e+17, 1.304322800397007e+17, 1.304322800470445e+17, 1.304322800547008e+17, 1.304322800620444e+17, 1.304322800693883e+17, 1.304322800765757e+17, 1.304322800840758e+17, 1.304322800912632e+17, 1.30432280098607e+17, 1.304322801064195e+17, 1.304322801142319e+17, 1.304322801215757e+17, 1.304322801290758e+17, 1.304322801362632e+17, 1.304322801437633e+17, 1.304322801512632e+17, 1.30432280158607e+17, 1.304322801662633e+17, 1.30432280173607e+17, 1.304322801807945e+17, 1.304322801886071e+17, 1.304322801957944e+17, 1.304322802031383e+17, 1.304322802109508e+17, 1.304322802182945e+17, 1.304322802256383e+17, 1.304322802331383e+17, 1.30432280240482e+17, 1.304322802478257e+17, 1.304322802556383e+17, 1.30432280262982e+17, 1.304322802703258e+17, 1.304322802778258e+17, 1.304322802851695e+17, 1.304322802925133e+17, 1.304322803003258e+17, 1.304322803076695e+17, 1.304322803150132e+17, 1.304322803225133e+17, 1.30432280329857e+17, 1.304322803372008e+17, 1.304322803462633e+17, 1.304322803542319e+17, 1.304322803614195e+17, 1.304322803695444e+17, 1.30432280376732e+17, 1.304322803840756e+17, 1.304322803915758e+17, 1.304322803989196e+17, 1.304322804062633e+17, 1.304322804140758e+17, 1.304322804212632e+17, 1.304322804286071e+17, 1.304322804359508e+17, 1.304322804432945e+17, 1.304322804506383e+17, 1.304322804579821e+17, 1.304322804659507e+17, 1.304322804731383e+17, 1.30432280480482e+17, 1.304322804876695e+17, 1.304322804953257e+17, 1.304322805025133e+17, 1.304322805100133e+17, 1.304322805176695e+17, 1.304322805251695e+17, 1.304322805325133e+17, 1.30432280539857e+17, 1.304322805472008e+17, 1.304322805545445e+17, 1.304322805625133e+17, 1.304322805697007e+17, 1.304322805770445e+17, 1.304322805848571e+17, 1.304322805922008e+17, 1.304322805995444e+17, 1.304322806072008e+17, 1.304322806147008e+17, 1.304322806220445e+17, 1.304322806293883e+17, 1.304322806365757e+17, 1.304322806439195e+17, 1.304322806511069e+17, 1.30432280658607e+17, 1.304322806659507e+17, 1.304322806731382e+17, 1.304322806804819e+17, 1.304322806878257e+17, 1.304322806956383e+17, 1.30432280702982e+17, 1.304322807106383e+17, 1.304322807179821e+17, 1.304322807253257e+17, 1.304322807328257e+17, 1.304322807401695e+17, 1.304322807473569e+17, 1.304322807548571e+17, 1.304322807625133e+17, 1.304322807697007e+17, 1.304322807770445e+17, 1.304322807843882e+17, 1.30432280791732e+17, 1.304322807990757e+17, 1.304322808064196e+17, 1.304322808142319e+17, 1.304322808228257e+17, 1.304322808307945e+17, 1.304322808384507e+17, 1.30432280846107e+17, 1.304322808534508e+17, 1.304322808607945e+17, 1.304322808681382e+17, 1.304322808756383e+17, 1.304322808832945e+17, 1.30432280890482e+17, 1.304322808978258e+17, 1.304322809051695e+17, 1.304322809128257e+17, 1.30432280919857e+17, 1.304322809272008e+17, 1.304322809345445e+17, 1.304322809422007e+17, 1.304322809495444e+17, 1.30432280956732e+17, 1.304322809645445e+17, 1.304322809718883e+17, 1.30432280979232e+17, 1.304322809868883e+17, 1.304322809942321e+17, 1.304322810015758e+17, 1.30432281009232e+17, 1.304322810165757e+17, 1.304322810239195e+17, 1.304322810312632e+17, 1.304322810387633e+17, 1.304322810459507e+17, 1.304322810532945e+17, 1.304322810611071e+17, 1.304322810684508e+17, 1.304322810757944e+17, 1.304322810834508e+17, 1.304322810906382e+17, 1.30432281097982e+17, 1.304322811053258e+17, 1.304322811128257e+17, 1.304322811201695e+17, 1.304322811273571e+17, 1.304322811350132e+17, 1.304322811425133e+17, 1.304322811500133e+17, 1.304322811573571e+17, 1.304322811648571e+17, 1.304322811722008e+17, 1.30432281179857e+17, 1.304322811872008e+17, 1.304322811945445e+17, 1.30432281202357e+17, 1.30432281209857e+17, 1.304322812172008e+17, 1.304322812247007e+17, 1.304322812320444e+17, 1.304322812393882e+17, 1.304322812467319e+17, 1.304322812540758e+17, 1.304322812615758e+17, 1.304322812690757e+17, 1.304322812764195e+17, 1.304322812837632e+17, 1.304322812920445e+17, 1.304322813020444e+17, 1.304322813100133e+17, 1.304322813175133e+17, 1.304322813253258e+17, 1.304322813326696e+17, 1.304322813401695e+17, 1.304322813790757e+17, 1.304322813864195e+17, 1.304322813937632e+17, 1.304322814009508e+17, 1.304322814084508e+17, 1.304322814157946e+17, 1.30432281423607e+17, 1.304322814309508e+17, 1.304322814382945e+17, 1.304322814459507e+17, 1.304322814540758e+17, 1.304322814614195e+17, 1.304322814689194e+17, 1.304322814765757e+17, 1.304322814837632e+17, 1.304322814911071e+17, 1.304322814987633e+17, 1.304322815059507e+17, 1.304322815134508e+17, 1.304322815211071e+17, 1.304322815284508e+17, 1.304322815357944e+17, 1.304322815434508e+17, 1.304322815507945e+17, 1.304322815581382e+17, 1.304322815657946e+17, 1.304322815743882e+17, 1.304322815822008e+17, 1.304322815893883e+17, 1.304322815970445e+17, 1.304322816043882e+17, 1.304322816118883e+17, 1.30432281619232e+17, 1.304322816265757e+17, 1.304322816339196e+17, 1.304322816412634e+17, 1.304322816484508e+17, 1.304322816557946e+17, 1.304322816632945e+17, 1.304322816706382e+17, 1.30432281677982e+17, 1.304322816856383e+17, 1.304322816932945e+17, 1.304322817006382e+17, 1.304322817079821e+17, 1.304322817156383e+17, 1.304322817232945e+17, 1.30432281730482e+17, 1.304322817376695e+17, 1.304322817450132e+17, 1.304322817525133e+17, 1.304322817600132e+17, 1.304322817673569e+17, 1.304322817750132e+17, 1.30432281782357e+17, 1.304322817897007e+17, 1.304322817973571e+17, 1.30432281804857e+17, 1.304322818137633e+17, 1.304322818217321e+17, 1.304322818290757e+17, 1.304322818365757e+17, 1.304322818440758e+17, 1.304322818512632e+17, 1.30432281858607e+17, 1.304322818662633e+17, 1.304322818737632e+17, 1.304322818809508e+17, 1.30432281888607e+17, 1.30432281896107e+17, 1.30432281903607e+17, 1.304322819109508e+17, 1.304322819182945e+17, 1.304322819256383e+17, 1.304322819337632e+17, 1.304322819414195e+17, 1.304322819487633e+17, 1.304322819562632e+17, 1.304322819637633e+17, 1.304322819711071e+17, 1.304322819784508e+17, 1.304322819856383e+17, 1.304322819934508e+17, 1.304322820006382e+17, 1.30432282007982e+17, 1.304322820157944e+17, 1.304322820226696e+17, 1.304322820301695e+17, 1.304322820375132e+17, 1.304322820451695e+17, 1.304322820534508e+17, 1.304322820612632e+17, 1.30432282068607e+17, 1.30432282076107e+17, 1.30432282083607e+17, 1.304322820909508e+17, 1.304322820981382e+17, 1.304322821053258e+17, 1.304322821128257e+17, 1.304322821201695e+17, 1.304322821275132e+17, 1.30432282134857e+17, 1.304322821425133e+17, 1.30432282149857e+17, 1.304322821573569e+17, 1.304322821648571e+17, 1.304322821731382e+17, 1.304322821806383e+17, 1.304322821879821e+17, 1.30432282195482e+17, 1.304322822028257e+17, 1.304322822101695e+17, 1.304322822178258e+17, 1.304322822250134e+17, 1.304322822326694e+17, 1.304322822400132e+17, 1.304322822473569e+17, 1.304322822548571e+17, 1.304322822626696e+17, 1.304322822700133e+17, 1.304322822773571e+17, 1.304322822847008e+17, 1.304322822943884e+17, 1.30432282302357e+17, 1.304322823095446e+17, 1.304322823178257e+17, 1.30432282325482e+17, 1.304322823328257e+17, 1.304322823400133e+17, 1.304322823473571e+17, 1.304322823551695e+17, 1.304322823626694e+17, 1.304322823700132e+17, 1.304322823773569e+17, 1.304322823847008e+17, 1.30432282392357e+17, 1.304322823997007e+17, 1.304322824070445e+17, 1.304322824150132e+17, 1.30432282422982e+17, 1.304322824303258e+17, 1.304322824375132e+17, 1.304322824453257e+17, 1.304322824526694e+17, 1.304322824600133e+17, 1.304322824675133e+17, 1.304322824748571e+17, 1.30432282482357e+17, 1.30432282489857e+17, 1.304322824972008e+17, 1.304322825045445e+17, 1.304322825125133e+17, 1.30432282519857e+17, 1.304322825273569e+17, 1.304322825353257e+17, 1.30432282542982e+17, 1.304322825503258e+17, 1.304322825579821e+17, 1.304322825662632e+17, 1.30432282573607e+17, 1.304322825812632e+17, 1.30432282588607e+17, 1.30432282596107e+17, 1.304322826037632e+17, 1.304322826111069e+17, 1.304322826184507e+17, 1.30432282626107e+17, 1.304322826334508e+17, 1.304322826407945e+17, 1.304322826484508e+17, 1.304322826565757e+17, 1.304322826640756e+17, 1.304322826714195e+17, 1.304322826790757e+17, 1.304322826864195e+17, 1.304322826937632e+17, 1.304322827011069e+17, 1.304322827084507e+17, 1.304322827157946e+17, 1.304322827234508e+17, 1.304322827307945e+17, 1.304322827381382e+17, 1.304322827457944e+17, 1.304322827531383e+17, 1.304322827604819e+17, 1.304322827682945e+17, 1.30432282776732e+17, 1.304322827847008e+17, 1.304322827920444e+17, 1.30432282799857e+17, 1.304322828072008e+17, 1.304322828150132e+17, 1.30432282822357e+17, 1.304322828297007e+17, 1.304322828372006e+17, 1.304322828447008e+17, 1.304322828529819e+17, 1.304322828601695e+17, 1.304322828676695e+17, 1.304322828750132e+17, 1.30432282882357e+17, 1.304322828900132e+17, 1.304322828981382e+17, 1.304322829057944e+17, 1.304322829131382e+17, 1.304322829207945e+17, 1.304322829282944e+17, 1.304322829359507e+17, 1.304322829428257e+17, 1.304322829501695e+17, 1.304322829575132e+17, 1.304322829653257e+17, 1.304322829726694e+17, 1.304322829800132e+17, 1.304322829875133e+17, 1.304322829950132e+17, 1.30432283002357e+17, 1.30432283009857e+17, 1.304322830182945e+17, 1.304322830262633e+17, 1.304322830334508e+17, 1.304322830412632e+17, 1.304322830484508e+17, 1.304322830559507e+17, 1.304322830634508e+17, 1.304322830707945e+17, 1.304322830782945e+17, 1.304322830856383e+17, 1.304322830932945e+17, 1.304322831006382e+17, 1.30432283107982e+17, 1.30432283115482e+17, 1.304322831228257e+17, 1.304322831300132e+17, 1.304322831381384e+17, 1.304322831456383e+17, 1.304322831528257e+17, 1.304322831603256e+17, 1.304322831678258e+17, 1.304322831751695e+17, 1.304322831826696e+17, 1.304322831900133e+17, 1.304322831972008e+17, 1.304322832050132e+17, 1.304322832125133e+17, 1.30432283219857e+17, 1.304322832272008e+17, 1.304322832347008e+17, 1.304322832420445e+17, 1.304322832497007e+17, 1.304322832590757e+17, 1.304322832670445e+17, 1.304322832743882e+17, 1.304322832828257e+17, 1.304322832903258e+17, 1.304322832976695e+17, 1.304322833050132e+17, 1.304322833125133e+17, 1.304322833201695e+17, 1.304322833276695e+17, 1.304322833350132e+17, 1.30432283342357e+17, 1.304322833497007e+17, 1.304322833573571e+17, 1.304322833647008e+17, 1.304322833722008e+17, 1.304322833800133e+17, 1.304322833876695e+17, 1.304322833950132e+17, 1.304322834026694e+17, 1.304322834100132e+17, 1.304322834175133e+17, 1.304322834248571e+17, 1.304322834325133e+17, 1.30432283439857e+17, 1.304322834470445e+17, 1.30432283454857e+17, 1.30432283462357e+17, 1.304322834697007e+17, 1.304322834770446e+17, 1.304322834843884e+17, 1.304322834915758e+17, 1.304322834997007e+17, 1.304322835076695e+17, 1.304322835150132e+17, 1.30432283522982e+17, 1.304322835301695e+17, 1.304322835373571e+17, 1.30432283544857e+17, 1.304322835522007e+17, 1.304322835597007e+17, 1.304322835670445e+17, 1.304322835747007e+17, 1.304322835820444e+17, 1.304322835893883e+17, 1.304322835970445e+17, 1.304322836043882e+17, 1.30432283611732e+17, 1.30432283619857e+17, 1.304322836273569e+17, 1.304322836347007e+17, 1.304322836423571e+17, 1.304322836497007e+17, 1.304322836572008e+17, 1.304322836647008e+17, 1.304322836722008e+17, 1.304322836795444e+17, 1.304322836868883e+17, 1.304322836945445e+17, 1.304322837018883e+17, 1.30432283709232e+17, 1.30432283716732e+17, 1.304322837240758e+17, 1.304322837312632e+17, 1.30432283739857e+17, 1.304322837475132e+17, 1.30432283754857e+17, 1.304322837626696e+17, 1.304322837700133e+17, 1.304322837773571e+17, 1.304322837850132e+17, 1.304322837925133e+17, 1.304322838001695e+17, 1.304322838075133e+17, 1.304322838150132e+17, 1.304322838225132e+17, 1.304322838298569e+17, 1.304322838372008e+17, 1.30432283844857e+17, 1.304322838522007e+17, 1.304322838601695e+17, 1.304322838675132e+17, 1.304322838751695e+17, 1.304322838826694e+17, 1.304322838900132e+17, 1.30432283898607e+17, 1.304322839059508e+17, 1.304322839134508e+17, 1.304322839206382e+17, 1.304322839281382e+17, 1.30432283935482e+17, 1.304322839428257e+17, 1.30432283950482e+17, 1.304322839578257e+17, 1.304322839651695e+17, 1.304322839726694e+17, 1.304322839812632e+17, 1.304322839889194e+17, 1.304322839962632e+17, 1.304322840037633e+17, 1.304322840112632e+17, 1.304322840187633e+17, 1.30432284026107e+17, 1.304322840337633e+17, 1.304322840412632e+17, 1.30432284048607e+17, 1.304322840559507e+17, 1.304322840634508e+17, 1.304322840707945e+17, 1.304322840784508e+17, 1.304322840857946e+17, 1.30432284092982e+17, 1.304322841007945e+17, 1.304322841082945e+17, 1.304322841157944e+17, 1.304322841231382e+17, 1.304322841304819e+17, 1.304322841378257e+17, 1.304322841453258e+17, 1.304322841528257e+17, 1.304322841603256e+17, 1.304322841676695e+17, 1.304322841750132e+17, 1.304322841825133e+17, 1.304322841901695e+17, 1.304322841973569e+17, 1.304322842048571e+17, 1.30432284212357e+17, 1.30432284221732e+17, 1.304322842293883e+17, 1.30432284236732e+17, 1.304322842450132e+17, 1.304322842525133e+17, 1.304322842597007e+17, 1.304322842672008e+17, 1.304322842745445e+17, 1.304322842826696e+17, 1.304322842895444e+17, 1.304322842968882e+17, 1.304322843042319e+17, 1.304322843120444e+17, 1.304322843193882e+17, 1.304322843267319e+17, 1.304322843343884e+17, 1.304322843425132e+17, 1.304322843498569e+17, 1.304322843572008e+17, 1.304322843650132e+17, 1.304322843725133e+17, 1.304322843797007e+17, 1.304322843870445e+17, 1.304322843945445e+17, 1.304322844015757e+17, 1.304322844089196e+17, 1.304322844164195e+17, 1.304322844237632e+17, 1.304322844311069e+17, 1.304322844384507e+17, 1.30432284446107e+17, 1.304322844532946e+17, 1.304322844614195e+17, 1.304322844687633e+17, 1.30432284476107e+17, 1.304322844837633e+17, 1.304322844907944e+17, 1.304322844981382e+17, 1.30432284505482e+17, 1.304322845131383e+17, 1.304322845206382e+17, 1.304322845278257e+17, 1.304322845353258e+17, 1.304322845426696e+17, 1.30432284549857e+17, 1.304322845572008e+17, 1.304322845647008e+17, 1.304322845722007e+17, 1.304322845797009e+17, 1.304322845873569e+17, 1.304322845945445e+17, 1.304322846018883e+17, 1.304322846097007e+17, 1.30432284616732e+17, 1.304322846240758e+17, 1.304322846314195e+17, 1.304322846389196e+17, 1.304322846462633e+17, 1.304322846537633e+17, 1.304322846612632e+17, 1.30432284668607e+17, 1.304322846759507e+17, 1.304322846837632e+17, 1.304322846911069e+17, 1.304322846990757e+17, 1.304322847065757e+17, 1.304322847140758e+17, 1.30432284721732e+17, 1.304322847290757e+17, 1.304322847362632e+17, 1.304322847437633e+17, 1.304322847509508e+17, 1.304322847582945e+17, 1.304322847656383e+17, 1.304322847731383e+17, 1.30432284780482e+17, 1.304322847876695e+17, 1.30432284795482e+17, 1.304322848028257e+17, 1.304322848100133e+17, 1.30432284817982e+17, 1.304322848253257e+17, 1.304322848325133e+17, 1.304322848400132e+17, 1.304322848473569e+17, 1.304322848547007e+17, 1.304322848625133e+17, 1.304322848698569e+17, 1.304322848772006e+17, 1.304322848848571e+17, 1.30432284892357e+17, 1.304322848995444e+17, 1.304322849072008e+17, 1.304322849145445e+17, 1.304322849220444e+17, 1.304322849293883e+17, 1.304322849370445e+17, 1.304322849447008e+17, 1.304322849520445e+17, 1.304322849600133e+17, 1.304322849673571e+17, 1.30432284974857e+17, 1.30432284982357e+17, 1.304322849897007e+17, 1.304322849970446e+17, 1.304322850047007e+17, 1.304322850120444e+17, 1.304322850195446e+17, 1.304322850268883e+17, 1.304322850342321e+17, 1.304322850415758e+17, 1.304322850489196e+17, 1.30432285056732e+17, 1.304322850643882e+17, 1.304322850717321e+17, 1.30432285079232e+17, 1.304322850865757e+17, 1.304322850939195e+17, 1.304322851014195e+17, 1.304322851084507e+17, 1.304322851164195e+17, 1.304322851237632e+17, 1.304322851311069e+17, 1.304322851387633e+17, 1.30432285146107e+17, 1.304322851534508e+17, 1.304322851611071e+17, 1.30432285168607e+17, 1.304322851772008e+17, 1.304322851848571e+17, 1.30432285192357e+17, 1.304322852006383e+17, 1.304322852078258e+17, 1.304322852151695e+17, 1.304322852231383e+17, 1.304322852303258e+17, 1.304322852376695e+17, 1.304322852451695e+17, 1.304322852525133e+17, 1.30432285259857e+17, 1.304322852672008e+17, 1.30432285274857e+17, 1.30432285282357e+17, 1.304322852897007e+17, 1.304322852973571e+17, 1.304322853047007e+17, 1.304322853125133e+17, 1.304322853195444e+17, 1.304322853268883e+17, 1.304322853342321e+17, 1.30432285341732e+17, 1.304322853490757e+17, 1.304322853564195e+17, 1.304322853642321e+17, 1.304322853715757e+17, 1.304322853789196e+17, 1.304322853864196e+17, 1.304322853937633e+17, 1.304322854011071e+17, 1.304322854082945e+17, 1.304322854164195e+17, 1.304322854240758e+17, 1.304322854314195e+17, 1.304322854393883e+17, 1.30432285446732e+17, 1.304322854540758e+17, 1.30432285461732e+17, 1.304322854690758e+17, 1.304322854767319e+17, 1.304322854839195e+17, 1.304322854912632e+17, 1.30432285498607e+17, 1.304322855059507e+17, 1.304322855132945e+17, 1.304322855206382e+17, 1.304322855279821e+17, 1.304322855359507e+17, 1.304322855432945e+17, 1.304322855506382e+17, 1.304322855582945e+17, 1.30432285565482e+17, 1.304322855728257e+17, 1.304322855801695e+17, 1.304322855875133e+17, 1.304322855948571e+17, 1.30432285602357e+17, 1.304322856100133e+17, 1.304322856173571e+17, 1.30432285624857e+17, 1.304322856322007e+17, 1.304322856395444e+17, 1.304322856468882e+17, 1.304322856553257e+17, 1.30432285662982e+17, 1.304322856703258e+17, 1.304322856781382e+17, 1.304322856853258e+17, 1.304322856926696e+17, 1.304322857000133e+17, 1.304322857073571e+17, 1.30432285714857e+17, 1.304322857226694e+17, 1.30432285729857e+17, 1.304322857372008e+17, 1.304322857445445e+17, 1.304322857520444e+17, 1.304322857595446e+17, 1.304322857665756e+17, 1.304322857747008e+17, 1.304322857820445e+17, 1.304322857893883e+17, 1.304322857968882e+17, 1.304322858042319e+17, 1.304322858115757e+17, 1.30432285819232e+17, 1.304322858265757e+17, 1.304322858339195e+17, 1.304322858415757e+17, 1.304322858489196e+17, 1.304322858562633e+17},
			             {1.304322320979821e+17, 1.304322321070445e+17, 1.30432232116107e+17, 1.304322321251695e+17, 1.304322321432945e+17},
			             {1.304322322518883e+17, 1.304322322609508e+17, 1.304322322700133e+17, 1.304322322790757e+17, 1.304322322881382e+17, 1.304322322972008e+17, 1.304322323062633e+17, 1.30432232315482e+17, 1.304322323243882e+17, 1.304322323334508e+17, 1.304322323425132e+17},
			             {1.304322331573571e+17, 1.304322331664196e+17, 1.304322331753257e+17, 1.30432233220482e+17},
			             {1.304322337275132e+17, 1.304322337365757e+17, 1.304322337454821e+17, 1.304322337545445e+17, 1.304322337637632e+17, 1.304322337728257e+17},
			             {1.30432234533607e+17, 1.304322345426694e+17, 1.304322345518883e+17, 1.304322345607945e+17, 1.304322345879821e+17, 1.304322345970445e+17},
			             {1.304322339356383e+17, 1.304322339718883e+17},
			             {1.304322358004819e+17, 1.304322358095444e+17, 1.304322358276695e+17},
			             {1.304322542589194e+17, 1.30432254421732e+17},
			             {1.30432256195482e+17, 1.304322562045445e+17, 1.304322562317321e+17, 1.304322562407945e+17, 1.30432256249857e+17, 1.304322562589196e+17, 1.30432256267982e+17, 1.304322562770445e+17, 1.30432256286107e+17, 1.304322563040758e+17, 1.304322563131383e+17},
			             {1.304322687582945e+17, 1.304322687659507e+17, 1.30432268772982e+17, 1.304322687803258e+17, 1.304322688097007e+17, 1.304322688170445e+17, 1.304322688318883e+17, 1.30432268839232e+17, 1.304322688465757e+17, 1.304322688540758e+17, 1.304322688837632e+17, 1.304322688909508e+17, 1.304322688987633e+17, 1.30432268906107e+17, 1.304322689134508e+17},
			             {1.304322708312632e+17, 1.304322708678258e+17, 1.304322708751695e+17, 1.304322708825133e+17, 1.304322709048571e+17, 1.304322709120445e+17, 1.304322709193883e+17, 1.304322709415757e+17},
			             {1.304322686489194e+17, 1.304322686562633e+17, 1.30432268663607e+17, 1.304322686709508e+17, 1.304322686781382e+17, 1.30432268685482e+17, 1.304322686928257e+17, 1.304322687000133e+17, 1.304322687073571e+17, 1.304322687147008e+17, 1.304322687220445e+17, 1.30432268772982e+17, 1.304322687803258e+17, 1.304322687875132e+17, 1.304322687951695e+17, 1.304322688025132e+17},
			             {1.304322688909508e+17, 1.304322688987633e+17, 1.30432268906107e+17, 1.304322689134508e+17, 1.304322689207945e+17, 1.304322689281382e+17, 1.304322689353258e+17, 1.304322689428257e+17, 1.304322689501695e+17, 1.304322689576695e+17, 1.304322690020445e+17, 1.30432269009232e+17, 1.304322690165757e+17, 1.304322690239196e+17, 1.304322690312634e+17},
			             {1.304322373207945e+17, 1.304322373478258e+17},
			             {1.30432261229232e+17, 1.304322612589196e+17},
			             {1.304322615689196e+17, 1.304322616059507e+17},
			             {1.30432261938607e+17, 1.304322620125132e+17},
			             {1.304322636815758e+17, 1.304322636890757e+17, 1.304322637111069e+17, 1.30432263718607e+17, 1.30432263741732e+17, 1.304322637490757e+17, 1.304322637564195e+17, 1.304322637637632e+17, 1.304322637712632e+17, 1.304322637931382e+17, 1.30432263800482e+17, 1.304322638079821e+17, 1.304322638153257e+17, 1.304322638226696e+17},
			             {1.304322647611071e+17, 1.304322649090757e+17},
			             {1.30432264938607e+17, 1.304322650420444e+17},
			             {1.304322649457944e+17, 1.304322650343884e+17},
			             {1.30432265286107e+17, 1.304322653598569e+17, 1.304322653672008e+17},
			             {1.304322639559507e+17, 1.304322640293882e+17},
			             {1.304322677665757e+17, 1.304322679070445e+17},
			             {1.30432267855482e+17, 1.304322679590757e+17},
			             {1.30432270270482e+17, 1.304322703228257e+17, 1.304322703301696e+17, 1.304322703376695e+17, 1.304322703453258e+17},
			             {1.30432275282357e+17, 1.304322753131383e+17, 1.304322753211069e+17, 1.304322753801695e+17},
			             {1.304322758456383e+17, 1.304322758531382e+17, 1.304322758603258e+17, 1.304322758681382e+17, 1.304322758753258e+17, 1.304322758826696e+17, 1.304322758900133e+17, 1.30432275898607e+17, 1.30432275913607e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}}, {{}, {}}, {{}, {}, {}}, {{}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}, {}}, {{}, {}}, {{}, {}}, {{}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
