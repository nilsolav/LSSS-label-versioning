netcdf mask {
	:date_created = "20200811T114915";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200811T114915";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 26;
			channels = 6;
			categories = 156;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  45.2, 32.9, 40.3, 49.1, 47.4, 49.1, 41.2, 51.7, 48.1, 49.2, 51.6, 45.7, 47.8, 49.9, 52.3, 46.4, 52.2, 55.9, 50.8, 49.7, 58.5, 55.5, 59.4, 53.6, 48.3, 51.9;
			max_depth =  50.0, 35.8, 44.2, 51.7, 52.1, 59.4, 48.3, 57.8, 55.2, 53.3, 54.6, 52.9, 50.7, 52.8, 56.0, 52.0, 55.9, 58.1, 55.7, 53.6, 60.3, 58.8, 61.4, 58.7, 58.3, 55.8;
			start_time = 131067418008401792, 131067417557308032, 131067418354339200, 131067418470745600, 131067430519964288, 131067430641526784, 131067427534495488, 131067427530276736, 131067427643714304, 131067427949182976, 131067422176683008, 131067423114339200, 131067419683870592, 131067424200901760, 131067425734964224, 131067426061839232, 131067431004495488, 131067431392464256, 131067431426683008, 131067431647620480, 131067431685745536, 131067424816214272, 131067432272464256, 131067432331995392, 131067432507776768, 131067432957151744;
			end_time = 131067418037620480, 131067417577464192, 131067418367620480, 131067418486995456, 131067430536214144, 131067430734339200, 131067427548089344, 131067427548089344, 131067427668558080, 131067427969964288, 131067422210120448, 131067423130901760, 131067419708401664, 131067424214026752, 131067425746995584, 131067426074339328, 131067431021995520, 131067431413245440, 131067431451526784, 131067431660120448, 131067431702464256, 131067424828401792, 131067432293870592, 131067432357151744, 131067432532151680, 131067432977933056;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21","Layer22","Layer23","Layer24","Layer25","Layer26";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63;
			mask_times = {1.310674180084018e+17, 1.310674180376205e+17},
			             {1.31067417557308e+17, 1.310674175774642e+17},
			             {1.310674183543392e+17, 1.310674183676205e+17},
			             {1.310674184707456e+17, 1.310674184869955e+17},
			             {1.310674305199643e+17, 1.310674305362141e+17},
			             {1.310674306415268e+17, 1.310674306459018e+17, 1.310674306499643e+17, 1.31067430654183e+17, 1.310674306584018e+17, 1.31067430662933e+17, 1.310674306671517e+17, 1.310674306712143e+17, 1.310674306752768e+17, 1.31067430679808e+17, 1.310674306838705e+17, 1.310674306879329e+17, 1.310674306921518e+17, 1.310674306962143e+17, 1.310674307002767e+17, 1.310674307048081e+17, 1.310674307088705e+17, 1.31067430712933e+17, 1.310674307169956e+17, 1.31067430721058e+17, 1.310674307259018e+17, 1.310674307302767e+17, 1.310674307343392e+17},
			             {1.310674275344955e+17, 1.310674275480893e+17},
			             {1.310674275302767e+17, 1.310674275480893e+17},
			             {1.310674276437143e+17, 1.310674276685581e+17},
			             {1.31067427949183e+17, 1.310674279699643e+17},
			             {1.31067422176683e+17, 1.310674221807456e+17, 1.310674221848079e+17, 1.310674221890267e+17, 1.310674221971517e+17, 1.310674222012142e+17, 1.31067422206058e+17, 1.310674222101204e+17},
			             {1.310674231143392e+17, 1.310674231309018e+17},
			             {1.310674196838706e+17, 1.310674197084017e+17},
			             {1.310674242009018e+17, 1.310674242140268e+17},
			             {1.310674257349642e+17, 1.310674257469956e+17},
			             {1.310674260618392e+17, 1.310674260743393e+17},
			             {1.310674310044955e+17, 1.310674310219955e+17},
			             {1.310674313924643e+17, 1.310674314132454e+17},
			             {1.31067431426683e+17, 1.310674314515268e+17},
			             {1.310674316476205e+17, 1.310674316601204e+17},
			             {1.310674316857455e+17, 1.310674317024643e+17},
			             {1.310674248162143e+17, 1.310674248284018e+17},
			             {1.310674322724643e+17, 1.31067432289183e+17, 1.310674322938706e+17},
			             {1.310674323319954e+17, 1.310674323571517e+17},
			             {1.310674325077768e+17, 1.310674325321517e+17},
			             {1.310674329571517e+17, 1.310674329779331e+17};
			mask_depths = {{45.2, 50.0}, {45.2, 50.0}}, {{32.9, 35.8}, {32.9, 35.8}}, {{40.3, 44.2}, {40.3, 44.2}}, {{49.1, 51.7}, {49.1, 51.7}}, {{47.4, 52.1}, {47.4, 52.1}}, {{49.1, 54.9}, {55.0, 55.3}, {55.4, 55.7}, {55.8, 56.0}, {56.1, 56.3}, {56.4, 56.7}, {56.8, 57.1}, {57.2, 57.3}, {57.4, 57.5}, {57.6, 57.8}, {49.1, 49.4, 57.9, 58.0}, {49.5, 50.1, 58.1, 58.4}, {50.2, 50.6}, {50.7, 51.1, 58.6, 58.7}, {51.2, 51.8, 58.8, 59.0}, {51.9, 52.1, 59.1, 59.2}, {52.2, 52.6, 59.3, 59.4}, {52.7, 52.9}, {53.0, 53.4}, {53.5, 54.4}, {54.5, 54.8}, {54.9, 55.2}, {55.3, 59.4}}, {{41.2, 48.3}, {41.2, 48.3}}, {{51.7, 57.8}, {51.7, 57.8}}, {{48.1, 55.2}, {48.1, 55.2}}, {{49.2, 53.3}, {49.2, 53.3}}, {{51.6, 54.5}, {54.4}, {54.4}, {54.5}, {54.5}, {54.6}, {54.5}, {51.6, 54.5}}, {{45.7, 52.9}, {45.7, 52.9}}, {{47.8, 50.7}, {47.8, 50.7}}, {{49.9, 52.8}, {49.9, 52.8}}, {{52.3, 56.0}, {52.3, 56.0}}, {{46.4, 52.0}, {46.4, 52.0}}, {{52.2, 55.9}, {52.2, 55.9}}, {{55.9, 58.1}, {55.9, 58.1}}, {{50.8, 55.7}, {50.8, 55.7}}, {{49.7, 53.6}, {49.7, 53.6}}, {{58.5, 60.3}, {58.5, 60.3}}, {{55.5, 58.8}, {55.5, 58.8}}, {{59.4, 61.4}, {61.4}, {59.4, 61.3}}, {{53.6, 58.7}, {53.6, 58.7}}, {{48.3, 58.3}, {48.3, 58.3}}, {{51.9, 55.8}, {51.9, 55.8}};
		}
	}
}
