netcdf mask {
	:date_created = "20200810T140900";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200810T140900";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 8;
			channels = 1;
			categories = 5;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  0.5, 10.4, 10.4, 10.4, 10.4, 41.6, 72.3,  0.0;
			max_depth =  10.4,  110.0,  109.0,  109.0,  109.0,   50.1,   80.3, 9999.0;
			start_time = 130590769912617216, 130590769912617216, 130590786276643968, 130590793269330176, 130590797170840320, 130590780599305600, 130590780696964608, 130590797178965504;
			end_time = 130590829941708032, 130590786276643968, 130590793269330176, 130590797170840320, 130590829941708032, 130590784354092928, 130590784696289408, 130590829941708032;
			region_id = 1, 2, 3, 4, 5, 6, 7, 8;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer1","Layer2","Layer1";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "";
			region_category_names = "0", "0", "0", "0", "0";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1, 2, 3, 4, 5;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "";
			region_channels = 1, 1, 1, 1, 1;
			mask_times = {1.305907699126172e+17, 1.305907699207424e+17, 1.305907699288677e+17, 1.305907699369929e+17, 1.305907699451181e+17, 1.305907699532433e+17, 1.305907699613684e+17, 1.305907699696499e+17, 1.305907699777751e+17, 1.305907699859003e+17, 1.305907699940256e+17, 1.305907700021508e+17, 1.30590770010276e+17, 1.305907700184013e+17, 1.305907700266828e+17, 1.305907700348079e+17, 1.305907700429332e+17, 1.305907700510583e+17, 1.305907700591836e+17, 1.305907700673088e+17, 1.30590770075434e+17, 1.305907700835592e+17, 1.305907700916844e+17, 1.305907700998095e+17, 1.305907701080911e+17, 1.305907701162163e+17, 1.305907701243415e+17, 1.305907701324667e+17, 1.305907701405919e+17, 1.305907701487172e+17, 1.305907701568424e+17, 1.305907701649676e+17, 1.305907701730929e+17, 1.30590770181218e+17, 1.305907701894995e+17, 1.305907701976248e+17, 1.3059077020575e+17, 1.305907702138752e+17, 1.305907702220004e+17, 1.305907702301256e+17, 1.305907702382508e+17, 1.305907702465322e+17, 1.305907702546575e+17, 1.305907702627827e+17, 1.305907702709079e+17, 1.305907702790331e+17, 1.305907702871583e+17, 1.305907702952835e+17, 1.305907703034088e+17, 1.30590770311534e+17, 1.305907703196591e+17, 1.305907703279406e+17, 1.305907703360658e+17, 1.305907703441911e+17, 1.305907703523164e+17, 1.305907703604416e+17, 1.305907703685668e+17, 1.30590770376692e+17, 1.305907703848172e+17, 1.305907703929423e+17, 1.305907704010675e+17, 1.30590770409349e+17, 1.305907704174742e+17, 1.305907704255995e+17, 1.305907704337247e+17, 1.3059077044185e+17, 1.30590770449975e+17, 1.305907704581004e+17, 1.305907704662255e+17, 1.30590770474507e+17, 1.305907704826322e+17, 1.305907704907575e+17, 1.305907704988827e+17, 1.305907705070079e+17, 1.305907705151332e+17, 1.305907705232584e+17, 1.305907705315398e+17, 1.30590770539665e+17, 1.305907705477902e+17, 1.305907705559154e+17, 1.305907705640406e+17, 1.305907705721658e+17, 1.305907705802909e+17, 1.305907705884163e+17, 1.305907705966977e+17, 1.305907706046668e+17, 1.305907706129482e+17, 1.305907706210734e+17, 1.305907706291986e+17, 1.305907706373238e+17, 1.305907706456052e+17, 1.305907706537306e+17, 1.305907706618557e+17, 1.305907706699809e+17, 1.305907706781062e+17, 1.305907706862314e+17, 1.305907706943566e+17, 1.305907707024818e+17, 1.305907707107633e+17, 1.305907707188886e+17, 1.305907707270136e+17, 1.305907707351388e+17, 1.305907707432641e+17, 1.305907707513893e+17, 1.305907707595145e+17, 1.305907707676398e+17, 1.30590770775765e+17, 1.305907707840465e+17, 1.305907707921716e+17, 1.305907708002968e+17, 1.305907708084221e+17, 1.305907708165473e+17, 1.305907708246725e+17, 1.305907708327978e+17, 1.30590770840923e+17, 1.305907708492045e+17, 1.305907708573297e+17, 1.305907708654548e+17, 1.3059077087358e+17, 1.305907708817052e+17, 1.305907708898304e+17, 1.305907708979557e+17, 1.305907709060809e+17, 1.305907709143624e+17, 1.305907709224876e+17, 1.305907709306127e+17, 1.30590770938738e+17, 1.305907709468632e+17, 1.305907709549884e+17, 1.305907709631137e+17, 1.305907709712389e+17, 1.305907709793641e+17, 1.305907709874893e+17, 1.305907709956145e+17, 1.305907710037398e+17, 1.305907710120212e+17, 1.305907710201464e+17, 1.305907710282716e+17, 1.305907710363968e+17, 1.30590771044522e+17, 1.305907710526473e+17, 1.305907710607725e+17, 1.305907710688977e+17, 1.305907710771791e+17, 1.305907710853044e+17, 1.305907710934296e+17, 1.305907711015548e+17, 1.3059077110968e+17, 1.305907711178053e+17, 1.305907711259305e+17, 1.30590771134212e+17, 1.305907711423372e+17, 1.305907711504623e+17, 1.305907711585876e+17, 1.305907711667128e+17, 1.305907711749943e+17, 1.305907711831195e+17, 1.305907711912447e+17, 1.305907711993699e+17, 1.30590771207495e+17, 1.305907712156202e+17, 1.305907712237455e+17, 1.305907712318707e+17, 1.305907712399959e+17, 1.305907712481212e+17, 1.305907712562464e+17, 1.305907712645279e+17, 1.305907712726531e+17, 1.305907712807784e+17, 1.305907712889036e+17, 1.305907712970287e+17, 1.305907713051539e+17, 1.305907713134354e+17, 1.305907713215607e+17, 1.305907713296859e+17, 1.305907713378111e+17, 1.305907713459363e+17, 1.305907713540614e+17, 1.305907713621866e+17, 1.305907713703118e+17, 1.305907713784371e+17, 1.305907713867185e+17, 1.305907713948438e+17, 1.305907714029691e+17, 1.305907714110943e+17, 1.305907714192195e+17, 1.305907714273446e+17, 1.3059077143547e+17, 1.305907714437513e+17, 1.305907714518766e+17, 1.305907714600018e+17, 1.30590771468127e+17, 1.305907714764084e+17, 1.305907714845338e+17, 1.305907714926589e+17, 1.305907715007841e+17, 1.305907715089093e+17, 1.305907715170345e+17, 1.305907715251597e+17, 1.30590771533285e+17, 1.305907715415665e+17, 1.305907715496916e+17, 1.305907715578168e+17, 1.30590771565942e+17, 1.305907715740673e+17, 1.305907715821925e+17, 1.305907715903177e+17, 1.305907715985992e+17, 1.305907716067244e+17, 1.305907716148497e+17, 1.305907716229748e+17, 1.305907716311e+17, 1.305907716392252e+17, 1.305907716473504e+17, 1.305907716554757e+17, 1.305907716637572e+17, 1.305907716718824e+17, 1.305907716800077e+17, 1.305907716881329e+17, 1.30590771696258e+17, 1.305907717045395e+17, 1.305907717126647e+17, 1.305907717207899e+17, 1.305907717289151e+17, 1.305907717370404e+17, 1.305907717453217e+17, 1.30590771753447e+17, 1.305907717615722e+17, 1.305907717696974e+17, 1.305907717778226e+17, 1.305907717859479e+17, 1.305907717940731e+17, 1.305907718021983e+17, 1.305907718104797e+17, 1.305907718186051e+17, 1.305907718267302e+17, 1.305907718348554e+17, 1.305907718431369e+17, 1.305907718512621e+17, 1.305907718593874e+17, 1.305907718675126e+17, 1.305907718756378e+17, 1.305907718837629e+17, 1.305907718918881e+17, 1.305907719000134e+17, 1.305907719082949e+17, 1.305907719164201e+17, 1.305907719245453e+17, 1.305907719326705e+17, 1.305907719407956e+17, 1.305907719489208e+17, 1.305907719570461e+17, 1.305907719651713e+17, 1.305907719734528e+17, 1.305907719815781e+17, 1.305907719897033e+17, 1.305907719978285e+17, 1.305907720059538e+17, 1.30590772014079e+17, 1.305907720222042e+17, 1.305907720303293e+17, 1.305907720386108e+17, 1.30590772046736e+17, 1.305907720548613e+17, 1.305907720629865e+17, 1.305907720711117e+17, 1.305907720792369e+17, 1.30590772087362e+17, 1.305907720954872e+17, 1.305907721037687e+17, 1.305907721118939e+17, 1.305907721200191e+17, 1.305907721281444e+17, 1.305907721362697e+17, 1.305907721443949e+17, 1.305907721525201e+17, 1.305907721606454e+17, 1.305907721687706e+17, 1.30590772177052e+17, 1.305907721851772e+17, 1.305907721933024e+17, 1.305907722014276e+17, 1.305907722097091e+17, 1.305907722178344e+17, 1.305907722259596e+17, 1.305907722340847e+17, 1.305907722422099e+17, 1.305907722503351e+17, 1.305907722584603e+17, 1.305907722667418e+17, 1.305907722748669e+17, 1.305907722829923e+17, 1.305907722911174e+17, 1.305907722992426e+17, 1.305907723073679e+17, 1.305907723154931e+17, 1.305907723236183e+17, 1.305907723317436e+17, 1.30590772340025e+17, 1.305907723481503e+17, 1.305907723562755e+17, 1.305907723644006e+17, 1.30590772372526e+17, 1.305907723806511e+17, 1.305907723887763e+17, 1.305907723969015e+17, 1.305907724050267e+17, 1.305907724133082e+17, 1.305907724214333e+17, 1.305907724295585e+17, 1.305907724376838e+17, 1.30590772445809e+17, 1.305907724539343e+17, 1.305907724620595e+17, 1.305907724701847e+17, 1.305907724784662e+17, 1.305907724865914e+17, 1.305907724947165e+17, 1.30590772502998e+17, 1.305907725111232e+17, 1.305907725192485e+17, 1.305907725273737e+17, 1.305907725354989e+17, 1.305907725436242e+17, 1.305907725517494e+17, 1.305907725600308e+17, 1.30590772568156e+17, 1.305907725762812e+17, 1.305907725844064e+17, 1.305907725925316e+17, 1.305907726006568e+17, 1.305907726087821e+17, 1.305907726169073e+17, 1.305907726251887e+17, 1.30590772633314e+17, 1.305907726414392e+17, 1.305907726495644e+17, 1.305907726576896e+17, 1.305907726658149e+17, 1.305907726739401e+17, 1.305907726820653e+17, 1.305907726903468e+17, 1.305907726984719e+17, 1.305907727065972e+17, 1.305907727147224e+17, 1.305907727228476e+17, 1.305907727309728e+17, 1.30590772739098e+17, 1.305907727472232e+17, 1.305907727553484e+17, 1.305907727634737e+17, 1.30590772771755e+17, 1.305907727798803e+17, 1.305907727880056e+17, 1.305907727961308e+17, 1.30590772804256e+17, 1.305907728125375e+17, 1.305907728205065e+17, 1.305907728287878e+17, 1.305907728369132e+17, 1.305907728450383e+17, 1.305907728531635e+17, 1.305907728612888e+17, 1.30590772869414e+17, 1.305907728775392e+17, 1.305907728856644e+17, 1.305907728937896e+17, 1.305907729019148e+17, 1.305907729101962e+17, 1.305907729183214e+17, 1.305907729264466e+17, 1.305907729345719e+17, 1.305907729428534e+17, 1.305907729509786e+17, 1.305907729591039e+17, 1.305907729672291e+17, 1.305907729753542e+17, 1.305907729834796e+17, 1.305907729916047e+17, 1.305907729997299e+17, 1.305907730078551e+17, 1.305907730159803e+17, 1.305907730241056e+17, 1.305907730323871e+17, 1.305907730405123e+17, 1.305907730486374e+17, 1.305907730567626e+17, 1.305907730648878e+17, 1.305907730730131e+17, 1.305907730811383e+17, 1.305907730894198e+17, 1.30590773097545e+17, 1.305907731056703e+17, 1.305907731137955e+17, 1.305907731219206e+17, 1.305907731300458e+17, 1.305907731381711e+17, 1.305907731464525e+17, 1.305907731545778e+17, 1.30590773162703e+17, 1.305907731708282e+17, 1.305907731789535e+17, 1.305907731870787e+17, 1.305907731952038e+17, 1.30590773203329e+17, 1.305907732114542e+17, 1.305907732195794e+17, 1.305907732278609e+17, 1.30590773235986e+17, 1.305907732441114e+17, 1.305907732522365e+17, 1.305907732603617e+17, 1.30590773268487e+17, 1.305907732766122e+17, 1.305907732847374e+17, 1.305907732930189e+17, 1.305907733011441e+17, 1.305907733092694e+17, 1.305907733173946e+17, 1.305907733255197e+17, 1.305907733336451e+17, 1.305907733417702e+17, 1.305907733500517e+17, 1.305907733580206e+17, 1.305907733663021e+17, 1.305907733744273e+17, 1.305907733825524e+17, 1.305907733906776e+17, 1.305907733988029e+17, 1.305907734070844e+17, 1.305907734150533e+17, 1.305907734231786e+17, 1.305907734314601e+17, 1.305907734395853e+17, 1.305907734477105e+17, 1.305907734558356e+17, 1.30590773463961e+17, 1.305907734722423e+17, 1.305907734803676e+17, 1.305907734884928e+17, 1.30590773496618e+17, 1.305907735047433e+17, 1.305907735128685e+17, 1.3059077352115e+17, 1.305907735292753e+17, 1.305907735374003e+17, 1.305907735455255e+17, 1.305907735536507e+17, 1.305907735617759e+17, 1.305907735700575e+17, 1.305907735781827e+17, 1.305907735863078e+17, 1.305907735944332e+17, 1.305907736027145e+17, 1.305907736108398e+17, 1.30590773618965e+17, 1.305907736270902e+17, 1.305907736352154e+17, 1.305907736433407e+17, 1.305907736514659e+17, 1.305907736595912e+17, 1.305907736678726e+17, 1.305907736759978e+17, 1.30590773684123e+17, 1.305907736922482e+17, 1.305907737003735e+17, 1.305907737084987e+17, 1.305907737166239e+17, 1.305907737247491e+17, 1.305907737328742e+17, 1.305907737411557e+17, 1.305907737492809e+17, 1.305907737574061e+17, 1.305907737655314e+17, 1.305907737736566e+17, 1.305907737817818e+17, 1.305907737900632e+17, 1.305907737981884e+17, 1.305907738063137e+17, 1.305907738144389e+17, 1.305907738225641e+17, 1.305907738306894e+17, 1.305907738388146e+17, 1.305907738469398e+17, 1.305907738550651e+17, 1.305907738633464e+17, 1.305907738714717e+17, 1.305907738795969e+17, 1.305907738877221e+17, 1.305907738960036e+17, 1.305907739041288e+17, 1.30590773912254e+17, 1.305907739203793e+17, 1.305907739285044e+17, 1.305907739366296e+17, 1.305907739447548e+17, 1.3059077395288e+17, 1.305907739611615e+17, 1.305907739692867e+17, 1.30590773977412e+17, 1.305907739855373e+17, 1.305907739936625e+17, 1.305907740017876e+17, 1.305907740099128e+17, 1.30590774018038e+17, 1.305907740263195e+17, 1.305907740344447e+17, 1.3059077404257e+17, 1.305907740506952e+17, 1.305907740588204e+17, 1.305907740669455e+17, 1.305907740750708e+17, 1.30590774083196e+17, 1.305907740914775e+17, 1.305907740996027e+17, 1.305907741077279e+17, 1.305907741158531e+17, 1.305907741241345e+17, 1.305907741322597e+17, 1.30590774140385e+17, 1.305907741485102e+17, 1.305907741566355e+17, 1.305907741647607e+17, 1.305907741728859e+17, 1.305907741811674e+17, 1.305907741892925e+17, 1.305907741974177e+17, 1.30590774205543e+17, 1.305907742136682e+17, 1.305907742217935e+17, 1.305907742300749e+17, 1.305907742382002e+17, 1.305907742463254e+17, 1.305907742544506e+17, 1.305907742625757e+17, 1.305907742707009e+17, 1.305907742788261e+17, 1.305907742869513e+17, 1.305907742950765e+17, 1.305907743032018e+17, 1.305907743113271e+17, 1.305907743196086e+17, 1.305907743277338e+17, 1.305907743358589e+17, 1.305907743439841e+17, 1.305907743521094e+17, 1.305907743602346e+17, 1.305907743683598e+17, 1.305907743766413e+17, 1.305907743847666e+17, 1.305907743928918e+17, 1.30590774401017e+17, 1.305907744091421e+17, 1.305907744172673e+17, 1.305907744253925e+17, 1.305907744335177e+17, 1.305907744417992e+17, 1.305907744499244e+17, 1.305907744580497e+17, 1.305907744661748e+17, 1.305907744743002e+17, 1.305907744825816e+17, 1.305907744907068e+17, 1.30590774498832e+17, 1.305907745069572e+17, 1.305907745150824e+17, 1.305907745232077e+17, 1.305907745313329e+17, 1.305907745394582e+17, 1.305907745475834e+17, 1.305907745557084e+17, 1.305907745638336e+17, 1.305907745719589e+17, 1.305907745800841e+17, 1.305907745883656e+17, 1.305907745964908e+17, 1.305907746046159e+17, 1.305907746127412e+17, 1.305907746208666e+17, 1.305907746289917e+17, 1.305907746371169e+17, 1.305907746453984e+17, 1.305907746535236e+17, 1.305907746616488e+17, 1.30590774669774e+17, 1.305907746778993e+17, 1.305907746861806e+17, 1.305907746943059e+17, 1.305907747024312e+17, 1.305907747105564e+17, 1.305907747186816e+17, 1.305907747268068e+17, 1.30590774734932e+17, 1.305907747430572e+17, 1.305907747511823e+17, 1.305907747593075e+17, 1.30590774767589e+17, 1.305907747757143e+17, 1.305907747838395e+17, 1.305907747919648e+17, 1.3059077480009e+17, 1.305907748082152e+17, 1.305907748163404e+17, 1.305907748244655e+17, 1.305907748325908e+17, 1.305907748408722e+17, 1.305907748489975e+17, 1.305907748571228e+17, 1.30590774865248e+17, 1.305907748733732e+17, 1.305907748814984e+17, 1.305907748896236e+17, 1.305907748977487e+17, 1.305907749060302e+17, 1.305907749141554e+17, 1.305907749222806e+17, 1.305907749304059e+17, 1.305907749385311e+17, 1.305907749466564e+17, 1.305907749549377e+17, 1.30590774963063e+17, 1.305907749711882e+17, 1.305907749793134e+17, 1.305907749875949e+17, 1.305907749957201e+17, 1.305907750038452e+17, 1.305907750119706e+17, 1.305907750200957e+17, 1.305907750282211e+17, 1.305907750363462e+17, 1.305907750446277e+17, 1.305907750527529e+17, 1.305907750608781e+17, 1.305907750690033e+17, 1.305907750771284e+17, 1.305907750852536e+17, 1.305907750933789e+17, 1.305907751015041e+17, 1.305907751096293e+17, 1.305907751177546e+17, 1.305907751258798e+17, 1.305907751341613e+17, 1.305907751422865e+17, 1.305907751504116e+17, 1.30590775158537e+17, 1.305907751666621e+17, 1.305907751747875e+17, 1.305907751829126e+17, 1.305907751911941e+17, 1.305907751993193e+17, 1.305907752074445e+17, 1.305907752155697e+17, 1.305907752236948e+17, 1.3059077523182e+17, 1.305907752399452e+17, 1.305907752480705e+17, 1.30590775256352e+17, 1.305907752644772e+17, 1.305907752726024e+17, 1.305907752807277e+17, 1.305907752888529e+17, 1.305907752971343e+17, 1.305907753052595e+17, 1.305907753133847e+17, 1.3059077532151e+17, 1.305907753296352e+17, 1.305907753377605e+17, 1.305907753458857e+17, 1.305907753541672e+17, 1.305907753622924e+17, 1.305907753704175e+17, 1.305907753785427e+17, 1.305907753866679e+17, 1.305907753947931e+17, 1.305907754029184e+17, 1.305907754111999e+17, 1.305907754193251e+17, 1.305907754274502e+17, 1.305907754355754e+17, 1.305907754437007e+17, 1.305907754518259e+17, 1.305907754599511e+17, 1.305907754680763e+17, 1.305907754762015e+17, 1.305907754844831e+17, 1.305907754926083e+17, 1.305907755007334e+17, 1.305907755088588e+17, 1.305907755169839e+17, 1.305907755251091e+17, 1.305907755332343e+17, 1.305907755413595e+17, 1.305907755494847e+17, 1.305907755577663e+17, 1.305907755658915e+17, 1.305907755740166e+17, 1.305907755821418e+17, 1.30590775590267e+17, 1.305907755983923e+17, 1.305907756065175e+17, 1.305907756146427e+17, 1.305907756229242e+17, 1.305907756310493e+17, 1.305907756391747e+17, 1.305907756472998e+17, 1.30590775655425e+17, 1.305907756635503e+17, 1.305907756716755e+17, 1.30590775679957e+17, 1.305907756880822e+17, 1.305907756962074e+17, 1.305907757043325e+17, 1.305907757124577e+17, 1.305907757207393e+17, 1.305907757288645e+17, 1.305907757369897e+17, 1.305907757451149e+17, 1.305907757532401e+17, 1.305907757613652e+17, 1.305907757694906e+17, 1.305907757776157e+17, 1.305907757858972e+17, 1.305907757940224e+17, 1.305907758021477e+17, 1.305907758102729e+17, 1.305907758183982e+17, 1.305907758265233e+17, 1.305907758346486e+17, 1.305907758427738e+17, 1.305907758508989e+17, 1.305907758591804e+17, 1.305907758673056e+17, 1.305907758754309e+17, 1.305907758835561e+17, 1.305907758916813e+17, 1.305907758998065e+17, 1.305907759079316e+17, 1.305907759160568e+17, 1.305907759241821e+17, 1.305907759323073e+17, 1.305907759404325e+17, 1.30590775948714e+17, 1.305907759568393e+17, 1.305907759649645e+17, 1.305907759730898e+17, 1.30590775981215e+17, 1.305907759893402e+17, 1.305907759974653e+17, 1.305907760055905e+17, 1.305907760137157e+17, 1.305907760218409e+17, 1.305907760301224e+17, 1.305907760382477e+17, 1.305907760463729e+17, 1.30590776054498e+17, 1.305907760626232e+17, 1.305907760707485e+17, 1.305907760788737e+17, 1.305907760869989e+17, 1.305907760951241e+17, 1.305907761034056e+17, 1.305907761115309e+17, 1.305907761196561e+17, 1.305907761277814e+17, 1.305907761359066e+17, 1.305907761440317e+17, 1.305907761521569e+17, 1.305907761602821e+17, 1.305907761684073e+17, 1.305907761765325e+17, 1.305907761846577e+17, 1.305907761929393e+17, 1.305907762010644e+17, 1.305907762091896e+17, 1.305907762173148e+17, 1.305907762254401e+17, 1.305907762335653e+17, 1.305907762416906e+17, 1.305907762498157e+17, 1.305907762580972e+17, 1.305907762662225e+17, 1.305907762743476e+17, 1.30590776282473e+17, 1.305907762905981e+17, 1.305907762987233e+17, 1.305907763068485e+17, 1.305907763149737e+17, 1.305907763230989e+17, 1.305907763312241e+17, 1.305907763395055e+17, 1.305907763476308e+17, 1.30590776355756e+17, 1.305907763638812e+17, 1.305907763720065e+17, 1.305907763801317e+17, 1.305907763882569e+17, 1.305907763963822e+17, 1.305907764046636e+17, 1.305907764127889e+17, 1.30590776420914e+17, 1.305907764290392e+17, 1.305907764371644e+17, 1.305907764452896e+17, 1.305907764534148e+17, 1.305907764616964e+17, 1.305907764698216e+17, 1.305907764779468e+17, 1.305907764860719e+17, 1.305907764941971e+17, 1.305907765023224e+17, 1.305907765104476e+17, 1.305907765185728e+17, 1.305907765266981e+17, 1.305907765349795e+17, 1.305907765431048e+17, 1.3059077655123e+17, 1.305907765593551e+17, 1.305907765674804e+17, 1.305907765756056e+17, 1.305907765837308e+17, 1.30590776591856e+17, 1.305907765999812e+17, 1.305907766081064e+17, 1.30590776616388e+17, 1.305907766245132e+17, 1.305907766326383e+17, 1.305907766407635e+17, 1.305907766488887e+17, 1.30590776657014e+17, 1.305907766651392e+17, 1.305907766734207e+17, 1.305907766815459e+17, 1.30590776689671e+17, 1.305907766979525e+17, 1.305907767060777e+17, 1.30590776714203e+17, 1.305907767223282e+17, 1.305907767304534e+17, 1.305907767385787e+17, 1.30590776746704e+17, 1.305907767549853e+17, 1.305907767631107e+17, 1.305907767712357e+17, 1.30590776779361e+17, 1.305907767874862e+17, 1.305907767956114e+17, 1.305907768037366e+17, 1.30590776812018e+17, 1.305907768201432e+17, 1.305907768282685e+17, 1.305907768363937e+17, 1.305907768446752e+17, 1.305907768528004e+17, 1.305907768609256e+17, 1.305907768690508e+17, 1.305907768771761e+17, 1.305907768853012e+17, 1.305907768934266e+17, 1.305907769015517e+17, 1.305907769096769e+17, 1.305907769179584e+17, 1.305907769260836e+17, 1.305907769342089e+17, 1.305907769423341e+17, 1.305907769504593e+17, 1.305907769585844e+17, 1.305907769668659e+17, 1.305907769749912e+17, 1.305907769831164e+17, 1.305907769912416e+17, 1.305907769993668e+17, 1.30590777007492e+17, 1.305907770156172e+17, 1.305907770238986e+17, 1.305907770320238e+17, 1.305907770401491e+17, 1.305907770482743e+17, 1.305907770563996e+17, 1.305907770645248e+17, 1.3059077707265e+17, 1.305907770807752e+17, 1.305907770889005e+17, 1.305907770970257e+17, 1.305907771051508e+17, 1.305907771134323e+17, 1.305907771215575e+17, 1.305907771296827e+17, 1.305907771378079e+17, 1.305907771459332e+17, 1.305907771540584e+17, 1.305907771621836e+17, 1.305907771703087e+17, 1.30590777178434e+17, 1.305907771867154e+17, 1.305907771948407e+17, 1.305907772029659e+17, 1.305907772110912e+17, 1.305907772192164e+17, 1.305907772274979e+17, 1.30590777235623e+17, 1.305907772437482e+17, 1.305907772518734e+17, 1.305907772599987e+17, 1.305907772681239e+17, 1.305907772764054e+17, 1.305907772845307e+17, 1.305907772926559e+17, 1.305907773007811e+17, 1.305907773089062e+17, 1.305907773170314e+17, 1.305907773251566e+17, 1.305907773334381e+17, 1.305907773415633e+17, 1.305907773496884e+17, 1.305907773578136e+17, 1.305907773659389e+17, 1.305907773740643e+17, 1.305907773821894e+17, 1.305907773903146e+17, 1.305907773984399e+17, 1.305907774065651e+17, 1.305907774146903e+17, 1.305907774229718e+17, 1.30590777431097e+17, 1.305907774392223e+17, 1.305907774473473e+17, 1.305907774554725e+17, 1.305907774635978e+17, 1.30590777471723e+17, 1.305907774798482e+17, 1.305907774879735e+17, 1.305907774962548e+17, 1.305907775043802e+17, 1.305907775125053e+17, 1.305907775206305e+17, 1.305907775287558e+17, 1.30590777536881e+17, 1.305907775450062e+17, 1.305907775531315e+17, 1.305907775612567e+17, 1.305907775695382e+17, 1.305907775776634e+17, 1.305907775857885e+17, 1.305907775939137e+17, 1.305907776020389e+17, 1.305907776101641e+17, 1.305907776182894e+17, 1.305907776264146e+17, 1.305907776345398e+17, 1.305907776428212e+17, 1.305907776509464e+17, 1.305907776590717e+17, 1.305907776671969e+17, 1.305907776753221e+17, 1.305907776834474e+17, 1.305907776917288e+17, 1.305907776998541e+17, 1.305907777079793e+17, 1.305907777161044e+17, 1.305907777242298e+17, 1.305907777323549e+17, 1.305907777404801e+17, 1.305907777486053e+17, 1.305907777567305e+17, 1.305907777648557e+17, 1.30590777772981e+17, 1.305907777811062e+17, 1.305907777892314e+17, 1.305907777975128e+17, 1.30590777805638e+17, 1.305907778137633e+17, 1.305907778218885e+17, 1.305907778300137e+17, 1.305907778382953e+17, 1.305907778462642e+17, 1.305907778543894e+17, 1.305907778626708e+17, 1.30590777870796e+17, 1.305907778789213e+17, 1.305907778870465e+17, 1.305907778951717e+17, 1.305907779032969e+17, 1.305907779114221e+17, 1.305907779195473e+17, 1.305907779276726e+17, 1.30590777935954e+17, 1.305907779440792e+17, 1.305907779522044e+17, 1.305907779604859e+17, 1.305907779686111e+17, 1.305907779767363e+17, 1.305907779848616e+17, 1.305907779929869e+17, 1.305907780011121e+17, 1.305907780092372e+17, 1.305907780173624e+17, 1.305907780254877e+17, 1.305907780336129e+17, 1.305907780418944e+17, 1.305907780500196e+17, 1.305907780581448e+17, 1.3059077806627e+17, 1.305907780743951e+17, 1.305907780825204e+17, 1.305907780906456e+17, 1.305907780987708e+17, 1.305907781068961e+17, 1.305907781150212e+17, 1.305907781231465e+17, 1.305907781312717e+17, 1.30590778139397e+17, 1.305907781475222e+17, 1.305907781558036e+17, 1.305907781639288e+17, 1.305907781720541e+17, 1.305907781801793e+17, 1.305907781884608e+17, 1.30590778196586e+17, 1.305907782047112e+17, 1.305907782128364e+17, 1.305907782209615e+17, 1.305907782290867e+17, 1.30590778237212e+17, 1.305907782453372e+17, 1.305907782534624e+17, 1.305907782615877e+17, 1.305907782697129e+17, 1.305907782779944e+17, 1.305907782861196e+17, 1.305907782942447e+17, 1.3059077830237e+17, 1.305907783104952e+17, 1.305907783186204e+17, 1.305907783267456e+17, 1.305907783350271e+17, 1.305907783431524e+17, 1.305907783512776e+17, 1.305907783594028e+17, 1.305907783675279e+17, 1.305907783756531e+17, 1.305907783837783e+17, 1.305907783919036e+17, 1.305907784000288e+17, 1.305907784083103e+17, 1.305907784164355e+17, 1.305907784245606e+17, 1.30590778432686e+17, 1.305907784408111e+17, 1.305907784489363e+17, 1.305907784570616e+17, 1.305907784651868e+17, 1.305907784734683e+17, 1.305907784815935e+17, 1.305907784897187e+17, 1.30590778497844e+17, 1.305907785059692e+17, 1.305907785140942e+17, 1.305907785222195e+17, 1.305907785303447e+17, 1.3059077853847e+17, 1.305907785465952e+17, 1.305907785547204e+17, 1.305907785630019e+17, 1.305907785709709e+17, 1.305907785792522e+17, 1.305907785873775e+17, 1.305907785955027e+17, 1.30590778603628e+17, 1.305907786117532e+17, 1.305907786198784e+17, 1.305907786280036e+17, 1.305907786362851e+17, 1.305907786444102e+17, 1.305907786525354e+17, 1.305907786606606e+17, 1.305907786687858e+17, 1.305907786769111e+17, 1.305907786850364e+17, 1.305907786931616e+17, 1.305907787012868e+17, 1.305907787095683e+17, 1.305907787176934e+17, 1.305907787258186e+17, 1.305907787339438e+17, 1.305907787420691e+17, 1.305907787501943e+17, 1.305907787584758e+17, 1.305907787666011e+17, 1.305907787747263e+17, 1.305907787828515e+17, 1.305907787909766e+17, 1.305907787992581e+17, 1.305907788073833e+17, 1.305907788155086e+17, 1.305907788236338e+17, 1.30590778831759e+17, 1.305907788398842e+17, 1.305907788480093e+17, 1.305907788561347e+17, 1.30590778864416e+17, 1.305907788725413e+17, 1.305907788806665e+17, 1.305907788887917e+17, 1.305907788969169e+17, 1.30590778905042e+17, 1.305907789131674e+17, 1.305907789212927e+17, 1.305907789294179e+17, 1.305907789376993e+17, 1.305907789458245e+17, 1.305907789539497e+17, 1.305907789620749e+17, 1.305907789702001e+17, 1.305907789784817e+17, 1.305907789866068e+17, 1.30590778994732e+17, 1.305907790028572e+17, 1.305907790109824e+17, 1.305907790192639e+17, 1.305907790272329e+17, 1.305907790355142e+17, 1.305907790434833e+17, 1.305907790517647e+17, 1.305907790598899e+17, 1.305907790680152e+17, 1.305907790761404e+17, 1.305907790842656e+17, 1.305907790923909e+17, 1.305907791005161e+17, 1.305907791086413e+17, 1.305907791167665e+17, 1.305907791248916e+17, 1.305907791330168e+17, 1.305907791412984e+17, 1.305907791494236e+17, 1.305907791575488e+17, 1.30590779165674e+17, 1.305907791737992e+17, 1.305907791819245e+17, 1.305907791900497e+17, 1.305907791981748e+17, 1.305907792063002e+17, 1.305907792145816e+17, 1.305907792227068e+17, 1.305907792308321e+17, 1.305907792389573e+17, 1.305907792470825e+17, 1.30590779255364e+17, 1.305907792634892e+17, 1.305907792716143e+17, 1.305907792797395e+17, 1.305907792878647e+17, 1.3059077929599e+17, 1.305907793041152e+17, 1.305907793122404e+17, 1.305907793203657e+17, 1.305907793284909e+17, 1.305907793367724e+17, 1.305907793448974e+17, 1.305907793530227e+17, 1.305907793611479e+17, 1.305907793692732e+17, 1.305907793773984e+17, 1.305907793856799e+17, 1.305907793938051e+17, 1.305907794019304e+17, 1.305907794100556e+17, 1.305907794181807e+17, 1.305907794263059e+17, 1.305907794344311e+17, 1.305907794427127e+17, 1.305907794508379e+17, 1.305907794589631e+17, 1.305907794670883e+17, 1.305907794752134e+17, 1.305907794833386e+17, 1.305907794914639e+17, 1.305907794995891e+17, 1.305907795078706e+17, 1.305907795159958e+17, 1.30590779524121e+17, 1.305907795322463e+17, 1.305907795403715e+17, 1.305907795484966e+17, 1.30590779556622e+17, 1.305907795647471e+17, 1.305907795728723e+17, 1.305907795809975e+17, 1.30590779589279e+17, 1.305907795974043e+17, 1.305907796055295e+17, 1.305907796136545e+17, 1.305907796217798e+17, 1.305907796300613e+17, 1.305907796381865e+17, 1.305907796463117e+17, 1.305907796544369e+17, 1.305907796625622e+17, 1.305907796706874e+17, 1.305907796788125e+17, 1.305907796870941e+17, 1.305907796952192e+17, 1.305907797033445e+17, 1.305907797114697e+17, 1.30590779719595e+17, 1.305907797277202e+17, 1.305907797360015e+17, 1.305907797441268e+17, 1.305907797522522e+17, 1.305907797603773e+17, 1.305907797685025e+17, 1.305907797766277e+17, 1.305907797847529e+17, 1.305907797928781e+17, 1.305907798010033e+17, 1.305907798092847e+17, 1.305907798174099e+17, 1.305907798255351e+17, 1.305907798336604e+17, 1.305907798417857e+17, 1.305907798499109e+17, 1.305907798580361e+17, 1.305907798663176e+17, 1.305907798742866e+17, 1.305907798825679e+17, 1.305907798906932e+17, 1.305907798988184e+17, 1.305907799069437e+17, 1.305907799152251e+17, 1.305907799233504e+17, 1.305907799314756e+17, 1.305907799396008e+17, 1.30590779947726e+17, 1.305907799558511e+17, 1.305907799639763e+17, 1.305907799722579e+17, 1.30590779980383e+17, 1.305907799885083e+17, 1.305907799966335e+17, 1.305907800047587e+17, 1.30590780012884e+17, 1.305907800210092e+17, 1.305907800291343e+17, 1.305907800372596e+17, 1.30590780045541e+17, 1.305907800536663e+17, 1.305907800617915e+17, 1.305907800699167e+17, 1.30590780078042e+17, 1.305907800861672e+17, 1.305907800942924e+17, 1.305907801025738e+17, 1.30590780110699e+17, 1.305907801188242e+17, 1.305907801269494e+17, 1.305907801350747e+17, 1.305907801431999e+17, 1.305907801513251e+17, 1.305907801594502e+17, 1.305907801675756e+17, 1.305907801758569e+17, 1.305907801839822e+17, 1.305907801921074e+17, 1.305907802002326e+17, 1.305907802083579e+17, 1.305907802164832e+17, 1.305907802246084e+17, 1.305907802327336e+17, 1.305907802408588e+17, 1.305907802489839e+17, 1.305907802571091e+17, 1.305907802653906e+17, 1.305907802735158e+17, 1.305907802816411e+17, 1.305907802897663e+17, 1.305907802978915e+17, 1.305907803060168e+17, 1.30590780314142e+17, 1.305907803224233e+17, 1.305907803305485e+17, 1.305907803386738e+17, 1.30590780346799e+17, 1.305907803550804e+17, 1.305907803632058e+17, 1.305907803713309e+17, 1.305907803794561e+17, 1.305907803875814e+17, 1.305907803955503e+17, 1.305907804038318e+17, 1.30590780411957e+17, 1.305907804200822e+17, 1.305907804283636e+17, 1.305907804364888e+17, 1.30590780444614e+17, 1.305907804527393e+17, 1.305907804608645e+17, 1.305907804689897e+17, 1.30590780477115e+17, 1.305907804852402e+17, 1.305907804935217e+17, 1.305907805016468e+17, 1.30590780509772e+17, 1.305907805178973e+17, 1.305907805260225e+17, 1.305907805341477e+17, 1.30590780542273e+17, 1.305907805503982e+17, 1.305907805586797e+17, 1.305907805668049e+17, 1.3059078057493e+17, 1.305907805830552e+17, 1.305907805911804e+17, 1.305907805993056e+17, 1.305907806074309e+17, 1.305907806155561e+17, 1.305907806236813e+17, 1.305907806318066e+17, 1.305907806400879e+17, 1.305907806482132e+17, 1.305907806563384e+17, 1.305907806644637e+17, 1.305907806725889e+17, 1.305907806807141e+17, 1.305907806888393e+17, 1.305907806969646e+17, 1.305907807050898e+17, 1.305907807133713e+17, 1.305907807214964e+17, 1.305907807296216e+17, 1.305907807377468e+17, 1.305907807458721e+17, 1.305907807541535e+17, 1.305907807622788e+17, 1.30590780770404e+17, 1.305907807785292e+17, 1.305907807866543e+17, 1.305907807947795e+17, 1.305907808029048e+17, 1.305907808111862e+17, 1.305907808193115e+17, 1.305907808272805e+17, 1.30590780835562e+17, 1.305907808436872e+17, 1.305907808518124e+17, 1.305907808599375e+17, 1.305907808680628e+17, 1.305907808763442e+17, 1.305907808844695e+17, 1.305907808925947e+17, 1.305907809007199e+17, 1.305907809088451e+17, 1.305907809169704e+17, 1.305907809250956e+17, 1.305907809332207e+17, 1.305907809413459e+17, 1.305907809496274e+17, 1.305907809577526e+17, 1.305907809658779e+17, 1.305907809740031e+17, 1.305907809821284e+17, 1.305907809902536e+17, 1.305907809983788e+17, 1.305907810065041e+17, 1.305907810146292e+17, 1.305907810229107e+17, 1.305907810310359e+17, 1.305907810391611e+17, 1.305907810472863e+17, 1.305907810554115e+17, 1.305907810635366e+17, 1.30590781071662e+17, 1.305907810797871e+17, 1.305907810880686e+17, 1.305907810961938e+17, 1.30590781104319e+17, 1.305907811124443e+17, 1.305907811205695e+17, 1.305907811286948e+17, 1.3059078113682e+17, 1.305907811449452e+17, 1.305907811532266e+17, 1.305907811613518e+17, 1.30590781169477e+17, 1.305907811776023e+17, 1.305907811857275e+17, 1.305907811938527e+17, 1.305907812019779e+17, 1.30590781210103e+17, 1.305907812183845e+17, 1.305907812265097e+17, 1.305907812346349e+17, 1.305907812427602e+17, 1.305907812508854e+17, 1.305907812591668e+17, 1.305907812671359e+17, 1.305907812752612e+17, 1.305907812833864e+17, 1.305907812916678e+17, 1.305907812996367e+17, 1.305907813079182e+17, 1.305907813160434e+17, 1.305907813241686e+17, 1.305907813322939e+17, 1.305907813405752e+17, 1.305907813485443e+17, 1.305907813568257e+17, 1.305907813649509e+17, 1.305907813730761e+17, 1.305907813812014e+17, 1.305907813893265e+17, 1.305907813974518e+17, 1.305907814057331e+17, 1.305907814138584e+17, 1.305907814219837e+17, 1.305907814301089e+17, 1.305907814382341e+17, 1.305907814463594e+17, 1.305907814546408e+17, 1.305907814627661e+17, 1.305907814708913e+17, 1.305907814790164e+17, 1.305907814871416e+17, 1.305907814952668e+17, 1.305907815033921e+17, 1.305907815116736e+17, 1.305907815197988e+17, 1.30590781527924e+17, 1.305907815360492e+17, 1.305907815441743e+17, 1.305907815522996e+17, 1.305907815604248e+17, 1.3059078156855e+17, 1.305907815766753e+17, 1.305907815849567e+17, 1.30590781593082e+17, 1.305907816012072e+17, 1.305907816093324e+17, 1.305907816174577e+17, 1.305907816255828e+17, 1.305907816338643e+17, 1.305907816419896e+17, 1.305907816501148e+17, 1.3059078165824e+17, 1.305907816663652e+17, 1.305907816744904e+17, 1.305907816826156e+17, 1.305907816907407e+17, 1.305907816988659e+17, 1.305907817071475e+17, 1.305907817152727e+17, 1.305907817233979e+17, 1.305907817315232e+17, 1.305907817396484e+17, 1.305907817477736e+17, 1.305907817558988e+17, 1.305907817641802e+17, 1.305907817723055e+17, 1.305907817804307e+17, 1.305907817885559e+17, 1.305907817966812e+17, 1.305907818048064e+17, 1.305907818129316e+17, 1.305907818210568e+17, 1.30590781829182e+17, 1.305907818373071e+17, 1.305907818455887e+17, 1.305907818537138e+17, 1.305907818618391e+17, 1.305907818699643e+17, 1.305907818780895e+17, 1.305907818862148e+17, 1.305907818943401e+17, 1.305907819024652e+17, 1.305907819107468e+17, 1.305907819188718e+17, 1.305907819269971e+17, 1.305907819351223e+17, 1.305907819432475e+17, 1.305907819513728e+17, 1.30590781959498e+17, 1.305907819676232e+17, 1.305907819759046e+17, 1.305907819840298e+17, 1.30590781992155e+17, 1.305907820002802e+17, 1.305907820084054e+17, 1.305907820165307e+17, 1.30590782024656e+17, 1.305907820329373e+17, 1.305907820410627e+17, 1.305907820491878e+17, 1.30590782057313e+17, 1.305907820654383e+17, 1.305907820737197e+17, 1.305907820816887e+17, 1.305907820899702e+17, 1.305907820980955e+17, 1.305907821062207e+17, 1.305907821143459e+17, 1.30590782122471e+17, 1.305907821305962e+17, 1.305907821388777e+17, 1.30590782147003e+17, 1.305907821551282e+17, 1.305907821632534e+17, 1.305907821713786e+17, 1.305907821795039e+17, 1.305907821876291e+17, 1.305907821959105e+17, 1.305907822040357e+17, 1.305907822121609e+17, 1.305907822202862e+17, 1.305907822284114e+17, 1.305907822365366e+17, 1.305907822446619e+17, 1.305907822527871e+17, 1.305907822609123e+17, 1.305907822691937e+17, 1.305907822773189e+17, 1.305907822854442e+17, 1.305907822935694e+17, 1.305907823016945e+17, 1.305907823099761e+17, 1.30590782317945e+17, 1.305907823262264e+17, 1.305907823343516e+17, 1.305907823424769e+17, 1.305907823507584e+17, 1.305907823588836e+17, 1.305907823670088e+17, 1.30590782375134e+17, 1.305907823832593e+17, 1.305907823913844e+17, 1.305907823995096e+17, 1.305907824076348e+17, 1.305907824159164e+17, 1.305907824240416e+17, 1.305907824321668e+17, 1.305907824402921e+17, 1.305907824484173e+17, 1.305907824565425e+17, 1.305907824646676e+17, 1.305907824729491e+17, 1.305907824810743e+17, 1.305907824891995e+17, 1.305907824974811e+17, 1.305907825056063e+17, 1.305907825137315e+17, 1.305907825218566e+17, 1.305907825299818e+17, 1.30590782538107e+17, 1.305907825462323e+17, 1.305907825543575e+17, 1.30590782562639e+17, 1.305907825707642e+17, 1.305907825788895e+17, 1.305907825870147e+17, 1.305907825951398e+17, 1.305907826032652e+17, 1.305907826113903e+17, 1.305907826195155e+17, 1.305907826276407e+17, 1.305907826359223e+17, 1.305907826440475e+17, 1.305907826521727e+17, 1.305907826602979e+17, 1.30590782668423e+17, 1.305907826765482e+17, 1.305907826846735e+17, 1.305907826927987e+17, 1.305907827010802e+17, 1.305907827092054e+17, 1.305907827173306e+17, 1.305907827254559e+17, 1.305907827335811e+17, 1.305907827417064e+17, 1.305907827498316e+17, 1.305907827579567e+17, 1.305907827660819e+17, 1.305907827742071e+17, 1.305907827824886e+17, 1.305907827906138e+17, 1.305907827987391e+17, 1.305907828068643e+17, 1.305907828149894e+17, 1.305907828231146e+17, 1.305907828312399e+17, 1.305907828393651e+17, 1.305907828474903e+17, 1.305907828557718e+17, 1.305907828638971e+17, 1.305907828720223e+17, 1.305907828801475e+17, 1.305907828882728e+17, 1.30590782896398e+17, 1.305907829045231e+17, 1.305907829126483e+17, 1.305907829207735e+17, 1.30590782929055e+17, 1.305907829371802e+17, 1.305907829453053e+17, 1.305907829534307e+17, 1.305907829615558e+17, 1.30590782969681e+17, 1.305907829778063e+17, 1.305907829859315e+17, 1.30590782994213e+17, 1.305907830023382e+17, 1.305907830104635e+17, 1.305907830187448e+17, 1.305907830268701e+17, 1.305907830349953e+17, 1.305907830431205e+17, 1.305907830512458e+17, 1.30590783059371e+17, 1.305907830674962e+17, 1.305907830756214e+17, 1.305907830837466e+17, 1.305907830920282e+17, 1.305907831001533e+17, 1.305907831082785e+17, 1.305907831164037e+17, 1.305907831245289e+17, 1.305907831326542e+17, 1.305907831407794e+17, 1.305907831489046e+17, 1.305907831570299e+17, 1.305907831651551e+17, 1.305907831734365e+17, 1.305907831815617e+17, 1.30590783189687e+17, 1.305907831978122e+17, 1.305907832059374e+17, 1.305907832140626e+17, 1.305907832221878e+17, 1.30590783230313e+17, 1.305907832384381e+17, 1.305907832467197e+17, 1.305907832546886e+17, 1.305907832629701e+17, 1.305907832710953e+17, 1.305907832792205e+17, 1.305907832873458e+17, 1.30590783295471e+17, 1.305907833035963e+17, 1.305907833117215e+17, 1.305907833200029e+17, 1.305907833281281e+17, 1.305907833362534e+17, 1.305907833443786e+17, 1.305907833525038e+17, 1.30590783360629e+17, 1.305907833687542e+17, 1.305907833768794e+17, 1.305907833851608e+17, 1.30590783393286e+17, 1.305907834014113e+17, 1.305907834095365e+17, 1.305907834176617e+17, 1.30590783425787e+17, 1.305907834339122e+17, 1.305907834421937e+17, 1.305907834503188e+17, 1.305907834584442e+17, 1.305907834665693e+17, 1.305907834746945e+17, 1.305907834828197e+17, 1.30590783490945e+17, 1.305907834990702e+17, 1.305907835071954e+17, 1.305907835154769e+17, 1.30590783523602e+17, 1.305907835317272e+17, 1.305907835398525e+17, 1.305907835479776e+17, 1.305907835561029e+17, 1.305907835642282e+17, 1.305907835723534e+17, 1.305907835806349e+17, 1.305907835887601e+17, 1.305907835968852e+17, 1.305907836050106e+17, 1.305907836131357e+17, 1.305907836212609e+17, 1.305907836293862e+17, 1.305907836375114e+17, 1.305907836456365e+17, 1.305907836537618e+17, 1.305907836620433e+17, 1.305907836701684e+17, 1.305907836782936e+17, 1.305907836864188e+17, 1.305907836945441e+17, 1.305907837026693e+17, 1.305907837107945e+17, 1.305907837189198e+17, 1.30590783727045e+17, 1.305907837351702e+17, 1.305907837432955e+17, 1.305907837514207e+17, 1.305907837597021e+17, 1.305907837678273e+17, 1.305907837759525e+17, 1.305907837840777e+17, 1.305907837922029e+17, 1.305907838003281e+17, 1.305907838084534e+17, 1.305907838165786e+17, 1.305907838247039e+17, 1.305907838328291e+17, 1.305907838411105e+17, 1.305907838492357e+17, 1.305907838573609e+17, 1.305907838654861e+17, 1.305907838736114e+17, 1.305907838817367e+17, 1.30590783890018e+17, 1.305907838979871e+17, 1.305907839062685e+17, 1.305907839143937e+17, 1.305907839225189e+17, 1.305907839306441e+17, 1.305907839387693e+17, 1.305907839468946e+17, 1.305907839550198e+17, 1.305907839633012e+17, 1.305907839714264e+17, 1.305907839795516e+17, 1.305907839876769e+17, 1.305907839958021e+17, 1.305907840039273e+17, 1.305907840120526e+17, 1.305907840203341e+17, 1.305907840284593e+17, 1.305907840365846e+17, 1.305907840447098e+17, 1.305907840528349e+17, 1.305907840609601e+17, 1.305907840692416e+17, 1.305907840773669e+17, 1.305907840854921e+17, 1.305907840936172e+17, 1.305907841017425e+17, 1.305907841098676e+17, 1.305907841179928e+17, 1.305907841261181e+17, 1.305907841342433e+17, 1.305907841425248e+17, 1.3059078415065e+17, 1.305907841587752e+17, 1.305907841669005e+17, 1.305907841750257e+17, 1.305907841831508e+17, 1.305907841912762e+17, 1.305907841994013e+17, 1.305907842075265e+17, 1.30590784215808e+17, 1.305907842239332e+17, 1.305907842320584e+17, 1.305907842401836e+17, 1.305907842484652e+17, 1.30590784256434e+17, 1.305907842645594e+17, 1.305907842726845e+17, 1.305907842808097e+17, 1.305907842889349e+17, 1.305907842972164e+17, 1.305907843053416e+17, 1.305907843134668e+17, 1.305907843215921e+17, 1.305907843297172e+17, 1.305907843378426e+17, 1.305907843459677e+17, 1.305907843540929e+17, 1.305907843622181e+17, 1.305907843704996e+17, 1.305907843786248e+17, 1.3059078438675e+17, 1.305907843948753e+17, 1.305907844030004e+17, 1.305907844111256e+17, 1.305907844192509e+17, 1.305907844273761e+17, 1.305907844355013e+17, 1.305907844437828e+17, 1.305907844519081e+17, 1.305907844600333e+17, 1.305907844681585e+17, 1.305907844762838e+17, 1.30590784484409e+17, 1.305907844925341e+17, 1.305907845006593e+17, 1.305907845087845e+17, 1.30590784517066e+17, 1.305907845251912e+17, 1.305907845333165e+17, 1.305907845414417e+17, 1.305907845495668e+17, 1.30590784557692e+17, 1.305907845658172e+17, 1.305907845739425e+17, 1.305907845820678e+17, 1.30590784590193e+17, 1.305907845984745e+17, 1.305907846065997e+17, 1.305907846147249e+17, 1.305907846228502e+17, 1.305907846309752e+17, 1.305907846392568e+17, 1.30590784647382e+17, 1.305907846555072e+17, 1.305907846636324e+17, 1.305907846717576e+17, 1.30590784680039e+17, 1.305907846881642e+17, 1.305907846962894e+17, 1.305907847044147e+17, 1.305907847125399e+17, 1.305907847206652e+17, 1.305907847287904e+17, 1.305907847369156e+17, 1.305907847450408e+17, 1.305907847533222e+17, 1.305907847614474e+17, 1.305907847695727e+17, 1.30590784777698e+17, 1.305907847858232e+17, 1.305907847939484e+17, 1.305907848020736e+17, 1.305907848101988e+17, 1.30590784818324e+17, 1.305907848264492e+17, 1.305907848347306e+17, 1.305907848428559e+17, 1.305907848509811e+17, 1.305907848591063e+17, 1.305907848672316e+17, 1.305907848753568e+17, 1.30590784883482e+17, 1.305907848916072e+17, 1.305907848997325e+17, 1.30590784908014e+17, 1.305907849161391e+17, 1.305907849242643e+17, 1.305907849323896e+17, 1.305907849405148e+17, 1.3059078494864e+17, 1.305907849567652e+17, 1.305907849650467e+17, 1.305907849731718e+17, 1.305907849812972e+17, 1.305907849894223e+17, 1.305907849975475e+17, 1.305907850056727e+17, 1.305907850137979e+17, 1.305907850219232e+17, 1.305907850300484e+17, 1.305907850381737e+17, 1.305907850464552e+17, 1.305907850545804e+17, 1.305907850627055e+17, 1.305907850708308e+17, 1.305907850789559e+17, 1.305907850870811e+17, 1.305907850952064e+17, 1.305907851033316e+17, 1.305907851114568e+17, 1.305907851197382e+17, 1.305907851278634e+17, 1.305907851359887e+17, 1.305907851442701e+17, 1.305907851523954e+17, 1.305907851605206e+17, 1.305907851686459e+17, 1.305907851767711e+17, 1.305907851847401e+17, 1.305907851930214e+17, 1.305907852011468e+17, 1.305907852092719e+17, 1.305907852173971e+17, 1.305907852255223e+17, 1.305907852338039e+17, 1.305907852419291e+17, 1.305907852500543e+17, 1.305907852581795e+17, 1.305907852663046e+17, 1.305907852744298e+17, 1.305907852827113e+17, 1.305907852908366e+17, 1.305907852989618e+17, 1.30590785307087e+17, 1.305907853152123e+17, 1.305907853233375e+17, 1.305907853314627e+17, 1.305907853397441e+17, 1.305907853478693e+17, 1.305907853559946e+17, 1.305907853641198e+17, 1.30590785372245e+17, 1.305907853803703e+17, 1.305907853884955e+17, 1.30590785396777e+17, 1.305907854047459e+17, 1.305907854130273e+17, 1.305907854211525e+17, 1.305907854292778e+17, 1.30590785437403e+17, 1.305907854455282e+17, 1.305907854536534e+17, 1.305907854619348e+17, 1.305907854700602e+17, 1.305907854781853e+17, 1.305907854863105e+17, 1.305907854944358e+17, 1.30590785502561e+17, 1.305907855108425e+17, 1.305907855189677e+17, 1.305907855270929e+17, 1.30590785535218e+17, 1.305907855433434e+17, 1.305907855514685e+17, 1.305907855595937e+17, 1.305907855677189e+17, 1.305907855760004e+17, 1.305907855841256e+17, 1.305907855922508e+17, 1.305907856003761e+17, 1.305907856085014e+17, 1.305907856166264e+17, 1.305907856247517e+17, 1.305907856330331e+17, 1.305907856411584e+17, 1.305907856492836e+17, 1.305907856574088e+17, 1.305907856655341e+17, 1.305907856736594e+17, 1.305907856819407e+17, 1.30590785690066e+17, 1.305907856981912e+17, 1.305907857063164e+17, 1.305907857145979e+17, 1.305907857227231e+17, 1.305907857308484e+17, 1.305907857389736e+17, 1.305907857470988e+17, 1.305907857552239e+17, 1.305907857633491e+17, 1.305907857716306e+17, 1.305907857797558e+17, 1.30590785787881e+17, 1.305907857960063e+17, 1.305907858041315e+17, 1.305907858122566e+17, 1.30590785820382e+17, 1.305907858285071e+17, 1.305907858367886e+17, 1.305907858449138e+17, 1.30590785853039e+17, 1.305907858611643e+17, 1.305907858692896e+17, 1.305907858775709e+17, 1.3059078588554e+17, 1.305907858938214e+17, 1.305907859019466e+17, 1.305907859100718e+17, 1.30590785918197e+17, 1.305907859263222e+17, 1.305907859346036e+17, 1.305907859427288e+17, 1.305907859508541e+17, 1.305907859589793e+17, 1.305907859671045e+17, 1.305907859752297e+17, 1.305907859835113e+17, 1.305907859916365e+17, 1.305907859997618e+17, 1.305907860078868e+17, 1.305907860160122e+17, 1.305907860241373e+17, 1.305907860322625e+17, 1.30590786040544e+17, 1.30590786048513e+17, 1.305907860567945e+17, 1.305907860649197e+17, 1.305907860730449e+17, 1.3059078608117e+17, 1.305907860894516e+17, 1.305907860975768e+17, 1.30590786105702e+17, 1.305907861138272e+17, 1.305907861219524e+17, 1.305907861300777e+17, 1.30590786138359e+17, 1.305907861464844e+17, 1.305907861546095e+17, 1.305907861627347e+17, 1.3059078617086e+17, 1.305907861789852e+17, 1.305907861871104e+17, 1.305907861952357e+17, 1.305907862033609e+17, 1.305907862114861e+17, 1.305907862196113e+17, 1.305907862277364e+17, 1.305907862358616e+17, 1.305907862441432e+17, 1.305907862522684e+17, 1.305907862603936e+17, 1.305907862685188e+17, 1.30590786276644e+17, 1.305907862847693e+17, 1.305907862930506e+17, 1.305907863011759e+17, 1.305907863093012e+17, 1.305907863174264e+17, 1.305907863255516e+17, 1.305907863336769e+17, 1.30590786341802e+17, 1.305907863499273e+17, 1.305907863580525e+17, 1.30590786366334e+17, 1.305907863744591e+17, 1.305907863825843e+17, 1.305907863908659e+17, 1.305907863989911e+17, 1.305907864071163e+17, 1.305907864152415e+17, 1.305907864233667e+17, 1.305907864314918e+17, 1.305907864396172e+17, 1.305907864478986e+17, 1.305907864560238e+17, 1.30590786464149e+17, 1.305907864722743e+17, 1.305907864803995e+17, 1.305907864885247e+17, 1.3059078649665e+17, 1.305907865047752e+17, 1.305907865129004e+17, 1.305907865210255e+17, 1.305907865293071e+17, 1.305907865374323e+17, 1.305907865455575e+17, 1.305907865536827e+17, 1.305907865618079e+17, 1.305907865699331e+17, 1.305907865780584e+17, 1.305907865861836e+17, 1.305907865943087e+17, 1.305907866025902e+17, 1.305907866107154e+17, 1.305907866188407e+17, 1.305907866269659e+17, 1.305907866350911e+17, 1.305907866432164e+17, 1.305907866513416e+17, 1.30590786659623e+17, 1.305907866677482e+17, 1.305907866758734e+17, 1.305907866839987e+17, 1.305907866921239e+17, 1.305907867004054e+17, 1.305907867085306e+17, 1.305907867166557e+17, 1.305907867247809e+17, 1.305907867329061e+17, 1.305907867410313e+17, 1.305907867491566e+17, 1.305907867572819e+17, 1.305907867654071e+17, 1.305907867735323e+17, 1.305907867816575e+17, 1.305907867899389e+17, 1.305907867980641e+17, 1.305907868061894e+17, 1.305907868143146e+17, 1.305907868224398e+17, 1.30590786830565e+17, 1.305907868386902e+17, 1.305907868469718e+17, 1.30590786855097e+17, 1.305907868632221e+17, 1.305907868713473e+17, 1.305907868794725e+17, 1.305907868875978e+17, 1.30590786895723e+17, 1.305907869038482e+17, 1.305907869119735e+17, 1.305907869200987e+17, 1.305907869282239e+17, 1.305907869363492e+17, 1.305907869444744e+17, 1.305907869525996e+17, 1.30590786960881e+17, 1.305907869690062e+17, 1.305907869771314e+17, 1.305907869852566e+17, 1.305907869933818e+17, 1.305907870015071e+17, 1.305907870096324e+17, 1.305907870177576e+17, 1.305907870258828e+17, 1.305907870341642e+17, 1.305907870422894e+17, 1.305907870504146e+17, 1.305907870586961e+17, 1.305907870668214e+17, 1.305907870749466e+17, 1.305907870830717e+17, 1.305907870911971e+17, 1.305907870993222e+17, 1.305907871074474e+17, 1.305907871155726e+17, 1.305907871238541e+17, 1.305907871319794e+17, 1.305907871401046e+17, 1.305907871482296e+17, 1.305907871563549e+17, 1.305907871644801e+17, 1.305907871726053e+17, 1.305907871807306e+17, 1.305907871888558e+17, 1.305907871971373e+17, 1.305907872052626e+17, 1.305907872133878e+17, 1.30590787221513e+17, 1.305907872296381e+17, 1.305907872377633e+17, 1.305907872458886e+17, 1.305907872540138e+17, 1.30590787262139e+17, 1.305907872704205e+17, 1.305907872785457e+17, 1.305907872866708e+17, 1.305907872947962e+17, 1.305907873029213e+17, 1.305907873110465e+17, 1.305907873191718e+17, 1.30590787327297e+17, 1.305907873355785e+17, 1.305907873437037e+17, 1.305907873518289e+17, 1.305907873599542e+17, 1.305907873680794e+17, 1.305907873762045e+17, 1.305907873843299e+17, 1.30590787392455e+17, 1.305907874005802e+17, 1.305907874088617e+17, 1.305907874169869e+17, 1.305907874251121e+17, 1.305907874332372e+17, 1.305907874413624e+17, 1.305907874494877e+17, 1.305907874576131e+17, 1.305907874658944e+17, 1.305907874740197e+17, 1.305907874821449e+17, 1.305907874902701e+17, 1.305907874983953e+17, 1.305907875065206e+17, 1.305907875146458e+17, 1.305907875227711e+17, 1.305907875308963e+17, 1.305907875391777e+17, 1.305907875473029e+17, 1.305907875554281e+17, 1.305907875635533e+17, 1.305907875716785e+17, 1.305907875799601e+17, 1.305907875880852e+17, 1.305907875962103e+17, 1.305907876043356e+17, 1.305907876124608e+17, 1.30590787620586e+17, 1.305907876288675e+17, 1.305907876368365e+17, 1.30590787645118e+17, 1.305907876532433e+17, 1.305907876613684e+17, 1.305907876694936e+17, 1.305907876776188e+17, 1.30590787685744e+17, 1.305907876938693e+17, 1.305907877019945e+17, 1.30590787710276e+17, 1.305907877184012e+17, 1.305907877265263e+17, 1.305907877346515e+17, 1.305907877427767e+17, 1.30590787750902e+17, 1.305907877590272e+17, 1.305907877671525e+17, 1.305907877752777e+17, 1.305907877835592e+17, 1.305907877916844e+17, 1.305907877998095e+17, 1.305907878079348e+17, 1.3059078781606e+17, 1.305907878241852e+17, 1.305907878323105e+17, 1.305907878404357e+17, 1.305907878485609e+17, 1.305907878568424e+17, 1.305907878649676e+17, 1.305907878730927e+17, 1.305907878812179e+17, 1.305907878893432e+17, 1.305907878974684e+17, 1.305907879055937e+17, 1.305907879137189e+17, 1.305907879218441e+17, 1.305907879299693e+17, 1.305907879380945e+17, 1.305907879463759e+17, 1.305907879545012e+17, 1.305907879626264e+17, 1.305907879707517e+17, 1.305907879788769e+17, 1.305907879870021e+17, 1.305907879952836e+17, 1.305907880034088e+17, 1.30590788011534e+17, 1.305907880196591e+17, 1.305907880277843e+17, 1.305907880360659e+17, 1.305907880441911e+17, 1.305907880523163e+17, 1.305907880604415e+17, 1.305907880685667e+17, 1.30590788076692e+17, 1.305907880848173e+17, 1.305907880929425e+17, 1.305907881010676e+17, 1.305907881093491e+17, 1.305907881174743e+17, 1.305907881255995e+17, 1.305907881337247e+17, 1.3059078814185e+17, 1.305907881499752e+17, 1.305907881582566e+17, 1.30590788166382e+17, 1.30590788174507e+17, 1.305907881826322e+17, 1.305907881907574e+17, 1.305907881988827e+17, 1.305907882070079e+17, 1.305907882152893e+17, 1.305907882234145e+17, 1.305907882315398e+17, 1.30590788239665e+17, 1.305907882477902e+17, 1.305907882559155e+17, 1.305907882641969e+17, 1.30590788272166e+17, 1.305907882802912e+17, 1.305907882884164e+17, 1.305907882966979e+17, 1.30590788304823e+17, 1.305907883129482e+17, 1.305907883210734e+17, 1.305907883291986e+17, 1.305907883373238e+17, 1.305907883454491e+17, 1.305907883535744e+17, 1.305907883618557e+17, 1.305907883699811e+17, 1.305907883781062e+17, 1.305907883863876e+17, 1.305907883943566e+17, 1.305907884026381e+17, 1.305907884107634e+17, 1.305907884188886e+17, 1.305907884270138e+17, 1.305907884351391e+17, 1.305907884432643e+17, 1.305907884513894e+17, 1.305907884595146e+17, 1.305907884676398e+17, 1.305907884759214e+17, 1.305907884840466e+17, 1.305907884921718e+17, 1.30590788500297e+17, 1.305907885084221e+17, 1.305907885165473e+17, 1.305907885246726e+17, 1.305907885329541e+17, 1.305907885410793e+17, 1.305907885492045e+17, 1.305907885573298e+17, 1.30590788565455e+17, 1.305907885735802e+17, 1.305907885817053e+17, 1.305907885898307e+17, 1.305907885981121e+17, 1.305907886062373e+17, 1.305907886143626e+17, 1.305907886224877e+17, 1.305907886306129e+17, 1.30590788638738e+17, 1.305907886468634e+17, 1.305907886549885e+17, 1.305907886631139e+17, 1.305907886713952e+17, 1.305907886795205e+17, 1.305907886876457e+17, 1.305907886957709e+17, 1.305907887038962e+17, 1.305907887120214e+17, 1.305907887201466e+17, 1.30590788728428e+17, 1.305907887365532e+17, 1.305907887446785e+17, 1.305907887528037e+17, 1.305907887609289e+17, 1.305907887690541e+17, 1.305907887771793e+17, 1.305907887854609e+17, 1.30590788793586e+17, 1.305907888017112e+17, 1.305907888098364e+17, 1.305907888179616e+17, 1.305907888260869e+17, 1.305907888343683e+17, 1.305907888424936e+17, 1.305907888506188e+17, 1.305907888587441e+17, 1.305907888668692e+17, 1.305907888749944e+17, 1.305907888831197e+17, 1.305907888912449e+17, 1.305907888993701e+17, 1.305907889076516e+17, 1.305907889157769e+17, 1.305907889239021e+17, 1.305907889320273e+17, 1.305907889401524e+17, 1.305907889482776e+17, 1.305907889564028e+17, 1.305907889646843e+17, 1.305907889728095e+17, 1.305907889809348e+17, 1.3059078898906e+17, 1.305907889971852e+17, 1.305907890053103e+17, 1.305907890134356e+17, 1.305907890215608e+17, 1.305907890296861e+17, 1.305907890379676e+17, 1.305907890460928e+17, 1.30590789054218e+17, 1.305907890623433e+17, 1.305907890704684e+17, 1.305907890785935e+17, 1.305907890867187e+17, 1.305907890948439e+17, 1.305907891029692e+17, 1.305907891112507e+17, 1.305907891193759e+17, 1.305907891275012e+17, 1.305907891356264e+17, 1.305907891437516e+17, 1.305907891518769e+17, 1.30590789160002e+17, 1.305907891681272e+17, 1.305907891762525e+17, 1.305907891843777e+17, 1.305907891926592e+17, 1.305907892007844e+17, 1.305907892089096e+17, 1.30590789217191e+17, 1.305907892253164e+17, 1.305907892334415e+17, 1.305907892415667e+17, 1.305907892496919e+17, 1.305907892578171e+17, 1.305907892659423e+17, 1.305907892740675e+17, 1.305907892821928e+17, 1.305907892904742e+17, 1.305907892985994e+17, 1.305907893067247e+17, 1.305907893148499e+17, 1.305907893229751e+17, 1.305907893311003e+17, 1.305907893392256e+17, 1.305907893475071e+17, 1.305907893556323e+17, 1.305907893637576e+17, 1.305907893718828e+17, 1.305907893800079e+17, 1.305907893882894e+17, 1.305907893964146e+17, 1.305907894045398e+17, 1.30590789412665e+17, 1.305907894207903e+17, 1.305907894289155e+17, 1.305907894370406e+17, 1.305907894451658e+17, 1.30590789453291e+17, 1.305907894614163e+17, 1.305907894696977e+17, 1.305907894776667e+17, 1.305907894859483e+17, 1.305907894940735e+17, 1.305907895021987e+17, 1.305907895104801e+17, 1.305907895186053e+17, 1.305907895267306e+17, 1.305907895348558e+17, 1.30590789542981e+17, 1.305907895511062e+17, 1.305907895592314e+17, 1.305907895673565e+17, 1.305907895754819e+17, 1.305907895837632e+17, 1.305907895918885e+17, 1.305907896000137e+17, 1.30590789608139e+17, 1.305907896162642e+17, 1.305907896243894e+17, 1.305907896325146e+17, 1.305907896406399e+17, 1.305907896489212e+17, 1.305907896570465e+17, 1.305907896651717e+17, 1.30590789673297e+17, 1.305907896814222e+17, 1.305907896895474e+17, 1.305907896976726e+17, 1.30590789705954e+17, 1.305907897140792e+17, 1.305907897222044e+17, 1.305907897303297e+17, 1.305907897384549e+17, 1.305907897465801e+17, 1.305907897547054e+17, 1.305907897628306e+17, 1.305907897709558e+17, 1.30590789779081e+17, 1.305907897872063e+17, 1.305907897954877e+17, 1.305907898036129e+17, 1.305907898117381e+17, 1.305907898198634e+17, 1.305907898279886e+17, 1.305907898361138e+17, 1.30590789844239e+17, 1.305907898523642e+17, 1.305907898604893e+17, 1.305907898686147e+17, 1.305907898767398e+17, 1.305907898850213e+17, 1.305907898931465e+17, 1.305907899012717e+17, 1.30590789909397e+17, 1.305907899175222e+17, 1.305907899256475e+17, 1.305907899337727e+17, 1.305907899418979e+17, 1.305907899501793e+17, 1.305907899583046e+17, 1.305907899664297e+17, 1.305907899745549e+17, 1.305907899826802e+17, 1.305907899908054e+17, 1.305907899990868e+17, 1.30590790007212e+17, 1.305907900153372e+17, 1.305907900234625e+17, 1.305907900317439e+17, 1.305907900398692e+17, 1.305907900479944e+17, 1.305907900561197e+17, 1.305907900642449e+17, 1.3059079007237e+17, 1.305907900804952e+17, 1.305907900886205e+17, 1.305907900969019e+17, 1.305907901050272e+17, 1.305907901131525e+17, 1.305907901212777e+17, 1.305907901294029e+17, 1.305907901375281e+17, 1.305907901458095e+17, 1.305907901539347e+17, 1.305907901620599e+17, 1.305907901701851e+17, 1.305907901784667e+17, 1.305907901865919e+17, 1.305907901947171e+17, 1.305907902028422e+17, 1.305907902109674e+17, 1.305907902190927e+17, 1.305907902272179e+17, 1.305907902353431e+17, 1.305907902434684e+17, 1.305907902515936e+17, 1.305907902597188e+17, 1.305907902680003e+17, 1.305907902759693e+17, 1.305907902842508e+17, 1.305907902922196e+17, 1.305907903005011e+17, 1.305907903086263e+17, 1.305907903167516e+17, 1.305907903248768e+17, 1.305907903331583e+17, 1.305907903412835e+17, 1.305907903492524e+17, 1.305907903573777e+17, 1.30590790365503e+17, 1.305907903737843e+17, 1.305907903819096e+17, 1.305907903900348e+17, 1.3059079039816e+17, 1.305907904062853e+17, 1.305907904144104e+17, 1.305907904225356e+17, 1.305907904306609e+17, 1.30590790438786e+17, 1.305907904470675e+17, 1.305907904551927e+17, 1.305907904633179e+17, 1.305907904714432e+17, 1.305907904797245e+17, 1.305907904878499e+17, 1.305907904958189e+17, 1.305907905039441e+17, 1.305907905122255e+17, 1.305907905201946e+17, 1.305907905284759e+17, 1.305907905364449e+17, 1.305907905447264e+17, 1.305907905528516e+17, 1.305907905609768e+17, 1.30590790569102e+17, 1.305907905772271e+17, 1.305907905853524e+17, 1.305907905934776e+17, 1.305907906017591e+17, 1.305907906098844e+17, 1.305907906180096e+17, 1.305907906261348e+17, 1.305907906342601e+17, 1.305907906423853e+17, 1.305907906506668e+17, 1.305907906587919e+17, 1.305907906669171e+17, 1.305907906750423e+17, 1.305907906831676e+17, 1.305907906912928e+17, 1.30590790699418e+17, 1.305907907075432e+17, 1.305907907156684e+17, 1.3059079072395e+17, 1.305907907319188e+17, 1.30590790740044e+17, 1.305907907481693e+17, 1.305907907562945e+17, 1.30590790764576e+17, 1.305907907727012e+17, 1.305907907808264e+17, 1.305907907889517e+17, 1.305907907970769e+17, 1.305907908053583e+17, 1.305907908134836e+17, 1.305907908216088e+17, 1.30590790829734e+17, 1.305907908378592e+17, 1.305907908459844e+17, 1.305907908542659e+17, 1.30590790862391e+17, 1.305907908705162e+17, 1.305907908786415e+17, 1.305907908867667e+17, 1.305907908948919e+17, 1.305907909030172e+17, 1.305907909111424e+17, 1.305907909192676e+17, 1.305907909275491e+17, 1.305907909356742e+17, 1.305907909437996e+17, 1.305907909519247e+17, 1.305907909600499e+17, 1.305907909681752e+17, 1.305907909763004e+17, 1.305907909844256e+17, 1.305907909927071e+17, 1.305907910008323e+17, 1.305907910089574e+17, 1.305907910170826e+17, 1.305907910252078e+17, 1.305907910333331e+17, 1.305907910414583e+17, 1.305907910495835e+17, 1.30590791057865e+17, 1.305907910659903e+17, 1.305907910741155e+17, 1.305907910822408e+17, 1.305907910903658e+17, 1.305907910984911e+17, 1.305907911066163e+17, 1.305907911147415e+17, 1.305907911230231e+17, 1.305907911311483e+17, 1.305907911392735e+17, 1.305907911473987e+17, 1.305907911555238e+17, 1.30590791163649e+17, 1.305907911719306e+17, 1.305907911800558e+17, 1.30590791188181e+17, 1.305907911963062e+17, 1.305907912044314e+17, 1.305907912125567e+17, 1.30590791220838e+17, 1.305907912289633e+17, 1.305907912370885e+17, 1.305907912452137e+17, 1.30590791253339e+17, 1.305907912614643e+17, 1.305907912695895e+17, 1.305907912777147e+17, 1.305907912859962e+17, 1.305907912941213e+17, 1.305907913022465e+17, 1.305907913103717e+17, 1.305907913184969e+17, 1.305907913266222e+17, 1.305907913347474e+17, 1.305907913430289e+17, 1.30590791351154e+17, 1.305907913592792e+17, 1.305907913674045e+17, 1.305907913755297e+17, 1.305907913836549e+17, 1.305907913917802e+17, 1.305907913999054e+17, 1.305907914080306e+17, 1.305907914163121e+17, 1.305907914244372e+17, 1.305907914325626e+17, 1.305907914406877e+17, 1.305907914488129e+17, 1.305907914569381e+17, 1.305907914650633e+17, 1.305907914733449e+17, 1.305907914814701e+17, 1.305907914895953e+17, 1.305907914977204e+17, 1.305907915058458e+17, 1.305907915139709e+17, 1.305907915220961e+17, 1.305907915303776e+17, 1.305907915385028e+17, 1.30590791546628e+17, 1.305907915547532e+17, 1.305907915628785e+17, 1.305907915710038e+17, 1.30590791579129e+17, 1.305907915872541e+17, 1.305907915955356e+17, 1.305907916036608e+17, 1.305907916117861e+17, 1.305907916199113e+17, 1.305907916280365e+17, 1.305907916361617e+17, 1.305907916442868e+17, 1.30590791652412e+17, 1.305907916606935e+17, 1.305907916688187e+17, 1.30590791676944e+17, 1.305907916850692e+17, 1.305907916931945e+17, 1.305907917013197e+17, 1.30590791709445e+17, 1.305907917175702e+17, 1.305907917256954e+17, 1.305907917338205e+17, 1.30590791742102e+17, 1.305907917502273e+17, 1.305907917583524e+17, 1.305907917664776e+17, 1.305907917746029e+17, 1.305907917827281e+17, 1.305907917910095e+17, 1.305907917991347e+17, 1.305907918072599e+17, 1.305907918153852e+17, 1.305907918235104e+17, 1.305907918316356e+17, 1.305907918397609e+17, 1.305907918478861e+17, 1.305907918560113e+17, 1.305907918642927e+17, 1.305907918724179e+17, 1.305907918805432e+17, 1.305907918886684e+17, 1.305907918967936e+17, 1.305907919050752e+17, 1.305907919132003e+17, 1.305907919211692e+17, 1.305907919294508e+17, 1.305907919375759e+17, 1.305907919457011e+17, 1.305907919538264e+17, 1.305907919619516e+17, 1.305907919702331e+17, 1.305907919783583e+17, 1.305907919864835e+17, 1.305907919946086e+17, 1.30590792002734e+17, 1.305907920110154e+17, 1.305907920191406e+17, 1.305907920272658e+17, 1.305907920353911e+17, 1.305907920435163e+17, 1.305907920516415e+17, 1.305907920597668e+17, 1.305907920680481e+17, 1.305907920761734e+17, 1.305907920842986e+17, 1.305907920924238e+17, 1.30590792100549e+17, 1.305907921088305e+17, 1.305907921169558e+17, 1.305907921250808e+17, 1.305907921332061e+17, 1.305907921413313e+17, 1.305907921494566e+17, 1.305907921575818e+17, 1.30590792165707e+17, 1.305907921738322e+17, 1.305907921821137e+17, 1.30590792190239e+17, 1.305907921983642e+17, 1.305907922064893e+17, 1.305907922146147e+17, 1.305907922227398e+17, 1.30590792230865e+17, 1.305907922391465e+17, 1.305907922472717e+17, 1.305907922553969e+17, 1.305907922635222e+17, 1.305907922716472e+17, 1.305907922797725e+17, 1.305907922878977e+17, 1.305907922960229e+17, 1.305907923043044e+17, 1.305907923124296e+17, 1.305907923205549e+17, 1.305907923286802e+17, 1.305907923368054e+17, 1.305907923449306e+17, 1.305907923530557e+17, 1.305907923611809e+17, 1.305907923693062e+17, 1.305907923774314e+17, 1.305907923855566e+17, 1.305907923936818e+17, 1.305907924019633e+17, 1.305907924100884e+17, 1.305907924182138e+17, 1.305907924263389e+17, 1.305907924344641e+17, 1.305907924425894e+17, 1.305907924507146e+17, 1.305907924588398e+17, 1.305907924671213e+17, 1.305907924752465e+17, 1.305907924833718e+17, 1.30590792491497e+17, 1.305907924996221e+17, 1.305907925077475e+17, 1.305907925158726e+17, 1.305907925239978e+17, 1.30590792532123e+17, 1.305907925404045e+17, 1.305907925485297e+17, 1.305907925566548e+17, 1.3059079256478e+17, 1.305907925729053e+17, 1.305907925810307e+17, 1.305907925891557e+17, 1.30590792597281e+17, 1.305907926055624e+17, 1.305907926136877e+17, 1.305907926218129e+17, 1.305907926299382e+17, 1.305907926380634e+17, 1.305907926461887e+17, 1.305907926543137e+17, 1.305907926624389e+17, 1.305907926705641e+17, 1.305907926788457e+17, 1.305907926869709e+17, 1.305907926950961e+17, 1.305907927032212e+17, 1.305907927113466e+17, 1.305907927196279e+17, 1.305907927277532e+17, 1.305907927357222e+17, 1.305907927440036e+17, 1.305907927521289e+17, 1.305907927602541e+17, 1.305907927683794e+17, 1.305907927765046e+17, 1.30590792784786e+17, 1.305907927929112e+17, 1.305907928010364e+17, 1.305907928091616e+17, 1.305907928213495e+17, 1.305907928336936e+17, 1.305907928457252e+17, 1.305907928538504e+17, 1.305907928621318e+17, 1.30590792870257e+17, 1.305907928783823e+17, 1.305907928863512e+17, 1.305907928946327e+17, 1.305907929027579e+17, 1.305907929108831e+17, 1.305907929190083e+17, 1.305907929271336e+17, 1.305907929352586e+17, 1.305907929433839e+17, 1.305907929516654e+17, 1.305907929597906e+17, 1.305907929679159e+17, 1.305907929760411e+17, 1.305907929841663e+17, 1.305907929922916e+17, 1.305907930005729e+17, 1.305907930086982e+17, 1.305907930168236e+17, 1.305907930249487e+17, 1.305907930330739e+17, 1.30590793041199e+17, 1.305907930493242e+17, 1.305907930574495e+17, 1.305907930657309e+17, 1.305907930738561e+17, 1.305907930819814e+17, 1.305907930901066e+17, 1.305907930982318e+17, 1.305907931063571e+17, 1.305907931144823e+17, 1.305907931226075e+17, 1.305907931307327e+17, 1.305907931390141e+17, 1.305907931471395e+17, 1.305907931552646e+17, 1.305907931633898e+17, 1.30590793171515e+17, 1.305907931796402e+17, 1.305907931877654e+17, 1.305907931958907e+17, 1.305907932041722e+17, 1.305907932122973e+17, 1.305907932204225e+17, 1.305907932285477e+17, 1.305907932368292e+17, 1.305907932449544e+17, 1.305907932530797e+17, 1.30590793261205e+17, 1.305907932693302e+17, 1.305907932774554e+17, 1.305907932857368e+17, 1.30590793293862e+17, 1.305907933019873e+17, 1.305907933101125e+17, 1.305907933182377e+17, 1.30590793326363e+17, 1.305907933344882e+17, 1.305907933426134e+17, 1.305907933507386e+17, 1.305907933588637e+17, 1.305907933671452e+17, 1.305907933752704e+17, 1.305907933833956e+17, 1.305907933915209e+17, 1.305907933996461e+17, 1.305907934077713e+17, 1.305907934158966e+17, 1.305907934240218e+17, 1.305907934323032e+17, 1.305907934404284e+17, 1.305907934485536e+17, 1.305907934566789e+17, 1.305907934649604e+17, 1.305907934730856e+17, 1.305907934812109e+17, 1.305907934893359e+17, 1.305907934974612e+17, 1.305907935055864e+17, 1.305907935138679e+17, 1.305907935219932e+17, 1.305907935301183e+17, 1.305907935382435e+17, 1.305907935463688e+17, 1.30590793554494e+17, 1.305907935626191e+17, 1.305907935707443e+17, 1.305907935788696e+17, 1.305907935869948e+17, 1.305907935952763e+17, 1.305907936034015e+17, 1.305907936115268e+17, 1.30590793619652e+17, 1.305907936277772e+17, 1.305907936359025e+17, 1.305907936440276e+17, 1.305907936521528e+17, 1.305907936604343e+17, 1.305907936685595e+17, 1.305907936766847e+17, 1.305907936848099e+17, 1.305907936930915e+17, 1.305907937010604e+17, 1.305907937093418e+17, 1.30590793717467e+17, 1.305907937255923e+17, 1.305907937337175e+17, 1.305907937418427e+17, 1.305907937501242e+17, 1.305907937582493e+17, 1.305907937663747e+17, 1.305907937744998e+17, 1.30590793782625e+17, 1.305907937907503e+17, 1.305907937988755e+17, 1.305907938070007e+17, 1.305907938152822e+17, 1.305907938234074e+17, 1.305907938315327e+17, 1.305907938396579e+17, 1.30590793847783e+17, 1.305907938559082e+17, 1.305907938640334e+17, 1.305907938721586e+17, 1.305907938804401e+17, 1.305907938885654e+17, 1.305907938966906e+17, 1.305907939048159e+17, 1.305907939129411e+17, 1.305907939210662e+17, 1.305907939291914e+17, 1.305907939373166e+17, 1.305907939454419e+17, 1.305907939537234e+17, 1.305907939618486e+17, 1.305907939699739e+17, 1.305907939780989e+17, 1.305907939862241e+17, 1.305907939943494e+17, 1.305907940024746e+17, 1.305907940105998e+17, 1.305907940187251e+17, 1.305907940268503e+17, 1.305907940351318e+17, 1.30590794043257e+17, 1.305907940513823e+17, 1.305907940595075e+17, 1.305907940676326e+17, 1.305907940757578e+17, 1.305907940838831e+17, 1.305907940920083e+17, 1.305907941001335e+17, 1.30590794108415e+17, 1.305907941165402e+17, 1.305907941246653e+17, 1.305907941327905e+17, 1.305907941409158e+17, 1.30590794149041e+17, 1.305907941571663e+17, 1.305907941652915e+17, 1.305907941734167e+17, 1.305907941816982e+17, 1.305907941898234e+17, 1.305907941979487e+17, 1.305907942060739e+17, 1.30590794214199e+17, 1.305907942223244e+17, 1.305907942304495e+17, 1.305907942385747e+17, 1.305907942466999e+17, 1.305907942548251e+17, 1.305907942629503e+17, 1.305907942712317e+17, 1.305907942793569e+17, 1.305907942874822e+17, 1.305907942956074e+17, 1.305907943037326e+17, 1.305907943118579e+17, 1.305907943199831e+17, 1.305907943281083e+17, 1.305907943362336e+17, 1.305907943443588e+17, 1.305907943526403e+17, 1.305907943607654e+17, 1.305907943688906e+17, 1.305907943770159e+17, 1.305907943851411e+17, 1.305907943932663e+17, 1.305907944013915e+17, 1.30590794409673e+17, 1.305907944177981e+17, 1.305907944259235e+17, 1.305907944340486e+17, 1.305907944423301e+17, 1.305907944504553e+17, 1.305907944585805e+17, 1.305907944667058e+17, 1.30590794474831e+17, 1.305907944829562e+17, 1.305907944912376e+17, 1.305907944993628e+17, 1.305907945074881e+17, 1.305907945156133e+17, 1.305907945237386e+17, 1.305907945318638e+17, 1.305907945401453e+17, 1.305907945482705e+17, 1.305907945563956e+17, 1.305907945645208e+17, 1.30590794572646e+17, 1.305907945807712e+17, 1.305907945888965e+17, 1.30590794597178e+17, 1.30590794605147e+17, 1.305907946134284e+17, 1.305907946215537e+17, 1.305907946296788e+17, 1.30590794637804e+17, 1.305907946460856e+17, 1.305907946542108e+17, 1.305907946621797e+17, 1.305907946704612e+17, 1.305907946785864e+17, 1.305907946867117e+17, 1.305907946948369e+17, 1.30590794702962e+17, 1.305907947110872e+17, 1.305907947192124e+17, 1.305907947273376e+17, 1.305907947354629e+17, 1.305907947435881e+17, 1.305907947517133e+17, 1.305907947598386e+17, 1.305907947679638e+17, 1.305907947762452e+17, 1.305907947843706e+17, 1.305907947924957e+17, 1.305907948006209e+17, 1.305907948087461e+17, 1.305907948168713e+17, 1.305907948249966e+17, 1.305907948331218e+17, 1.30590794841247e+17, 1.305907948493722e+17, 1.305907948576536e+17, 1.305907948657788e+17, 1.305907948739041e+17, 1.305907948820293e+17, 1.305907948901545e+17, 1.305907948982797e+17, 1.30590794906405e+17, 1.305907949145302e+17, 1.305907949228116e+17, 1.305907949309368e+17, 1.305907949390621e+17, 1.305907949473435e+17, 1.305907949554688e+17, 1.30590794963594e+17, 1.305907949717192e+17, 1.305907949798445e+17, 1.305907949879697e+17, 1.305907949960948e+17, 1.3059079500422e+17, 1.305907950123452e+17, 1.305907950204705e+17, 1.305907950285957e+17, 1.305907950368772e+17, 1.305907950450024e+17, 1.305907950531276e+17, 1.305907950612529e+17, 1.30590795069378e+17, 1.305907950775034e+17, 1.305907950857847e+17, 1.3059079509391e+17, 1.305907951020352e+17, 1.305907951101604e+17, 1.305907951182857e+17, 1.305907951264109e+17, 1.305907951345361e+17, 1.305907951428175e+17, 1.305907951509427e+17, 1.305907951590679e+17, 1.305907951671931e+17, 1.305907951753183e+17, 1.305907951834436e+17, 1.305907951915688e+17, 1.30590795199694e+17, 1.305907952078193e+17, 1.305907952159446e+17, 1.305907952242259e+17, 1.305907952323512e+17, 1.305907952404764e+17, 1.305907952486016e+17, 1.305907952567268e+17, 1.30590795264852e+17, 1.305907952729773e+17, 1.305907952811025e+17, 1.305907952893839e+17, 1.305907952975091e+17, 1.305907953056343e+17, 1.305907953137595e+17, 1.305907953218847e+17, 1.305907953301661e+17, 1.305907953381352e+17, 1.305907953464166e+17, 1.305907953545418e+17, 1.305907953626671e+17, 1.305907953707923e+17, 1.305907953789175e+17, 1.305907953870428e+17, 1.30590795395168e+17, 1.305907954034495e+17, 1.305907954115748e+17, 1.305907954196998e+17, 1.305907954278252e+17, 1.305907954359503e+17, 1.305907954440755e+17, 1.305907954522007e+17, 1.305907954604822e+17, 1.305907954686074e+17, 1.305907954767327e+17, 1.305907954848579e+17, 1.30590795492983e+17, 1.305907955011082e+17, 1.305907955092335e+17, 1.30590795517515e+17, 1.305907955256402e+17, 1.305907955337655e+17, 1.305907955418907e+17, 1.305907955500159e+17, 1.305907955581411e+17, 1.305907955662664e+17, 1.305907955743916e+17, 1.305907955825167e+17, 1.305907955906419e+17, 1.305907955989234e+17, 1.305907956070486e+17, 1.305907956151738e+17, 1.305907956232989e+17, 1.305907956314243e+17, 1.305907956395494e+17, 1.305907956476746e+17, 1.305907956557999e+17, 1.305907956639252e+17, 1.305907956720503e+17, 1.305907956801756e+17, 1.305907956883008e+17, 1.30590795696426e+17, 1.305907957047075e+17, 1.305907957128328e+17, 1.30590795720958e+17, 1.305907957290831e+17, 1.305907957372083e+17, 1.305907957453335e+17, 1.305907957534587e+17, 1.305907957617402e+17, 1.305907957698655e+17, 1.305907957779907e+17, 1.305907957861158e+17, 1.305907957942412e+17, 1.305907958023663e+17, 1.305907958104915e+17, 1.305907958186168e+17, 1.305907958268982e+17, 1.305907958350235e+17, 1.305907958431487e+17, 1.305907958512739e+17, 1.30590795859399e+17, 1.305907958675242e+17, 1.305907958756494e+17, 1.305907958837747e+17, 1.305907958918999e+17, 1.305907959000251e+17, 1.305907959083067e+17, 1.305907959164319e+17, 1.305907959245571e+17, 1.305907959326822e+17, 1.305907959408076e+17, 1.305907959489327e+17, 1.305907959570579e+17, 1.305907959651832e+17, 1.305907959734647e+17, 1.305907959815899e+17, 1.305907959897151e+17, 1.305907959978403e+17, 1.305907960059654e+17, 1.305907960140906e+17, 1.305907960222159e+17, 1.305907960303411e+17, 1.305907960386226e+17, 1.305907960467478e+17, 1.30590796054873e+17, 1.305907960629983e+17, 1.305907960712796e+17, 1.305907960794049e+17, 1.305907960875301e+17, 1.305907960956554e+17, 1.305907961037806e+17, 1.305907961119058e+17, 1.305907961200311e+17, 1.305907961283124e+17, 1.305907961364378e+17, 1.305907961445629e+17, 1.305907961526883e+17, 1.305907961608134e+17, 1.305907961689386e+17, 1.305907961770638e+17, 1.30590796185189e+17, 1.305907961934705e+17, 1.305907962015956e+17, 1.305907962097208e+17, 1.305907962178461e+17, 1.305907962259713e+17, 1.305907962340965e+17, 1.305907962422218e+17, 1.30590796250347e+17, 1.305907962584722e+17, 1.305907962667537e+17, 1.30590796274879e+17, 1.305907962830042e+17, 1.305907962911293e+17, 1.305907962992545e+17, 1.305907963073797e+17, 1.305907963155049e+17, 1.305907963237865e+17, 1.305907963319117e+17, 1.305907963400369e+17, 1.30590796348162e+17, 1.305907963564435e+17, 1.305907963645687e+17, 1.30590796372694e+17, 1.305907963808192e+17, 1.305907963889444e+17, 1.305907963970696e+17, 1.305907964051949e+17, 1.305907964133201e+17, 1.305907964214454e+17, 1.305907964297267e+17, 1.30590796437852e+17, 1.305907964459772e+17, 1.305907964541024e+17, 1.305907964622277e+17, 1.305907964701966e+17, 1.305907964784781e+17, 1.305907964866033e+17, 1.305907964947284e+17, 1.305907965030099e+17, 1.305907965111351e+17, 1.305907965192604e+17, 1.305907965273856e+17, 1.305907965355109e+17, 1.305907965436361e+17, 1.305907965517613e+17, 1.305907965598865e+17, 1.305907965680116e+17, 1.30590796576137e+17, 1.305907965842621e+17, 1.305907965923873e+17, 1.305907966005125e+17, 1.305907966087941e+17, 1.305907966169193e+17, 1.305907966250445e+17, 1.305907966331697e+17, 1.305907966412948e+17, 1.305907966494202e+17, 1.305907966577015e+17, 1.305907966658268e+17, 1.30590796673952e+17, 1.305907966820772e+17, 1.305907966902025e+17, 1.305907966983277e+17, 1.305907967064529e+17, 1.305907967147345e+17, 1.305907967228596e+17, 1.305907967309848e+17, 1.3059079673911e+17, 1.305907967472352e+17, 1.305907967553604e+17, 1.305907967634856e+17, 1.305907967716109e+17, 1.305907967798924e+17, 1.305907967880175e+17, 1.30590796796299e+17, 1.305907968044242e+17, 1.305907968125494e+17, 1.305907968206746e+17, 1.305907968287999e+17, 1.305907968369251e+17, 1.305907968450504e+17, 1.305907968533317e+17, 1.30590796861457e+17, 1.305907968695822e+17, 1.305907968777074e+17, 1.305907968858327e+17, 1.305907968939579e+17, 1.305907969020832e+17, 1.305907969102084e+17, 1.305907969184899e+17, 1.30590796926615e+17, 1.305907969347402e+17, 1.305907969428654e+17, 1.305907969509906e+17, 1.305907969591158e+17, 1.305907969672411e+17, 1.305907969753663e+17, 1.305907969834916e+17, 1.305907969916168e+17, 1.30590796999742e+17, 1.305907970078671e+17, 1.305907970159923e+17, 1.305907970242739e+17, 1.305907970323991e+17, 1.305907970405243e+17, 1.305907970486496e+17, 1.305907970567748e+17, 1.305907970649e+17, 1.305907970730252e+17, 1.305907970811503e+17, 1.305907970894318e+17, 1.30590797097557e+17, 1.305907971056822e+17, 1.305907971138075e+17, 1.305907971219327e+17, 1.305907971300579e+17, 1.305907971381832e+17, 1.305907971463084e+17, 1.305907971544335e+17, 1.305907971627151e+17, 1.305907971708403e+17, 1.305907971789655e+17, 1.305907971870907e+17, 1.305907971952159e+17, 1.305907972033411e+17, 1.305907972114662e+17, 1.305907972197478e+17, 1.30590797227873e+17, 1.305907972359982e+17, 1.305907972441234e+17, 1.305907972522486e+17, 1.3059079726053e+17, 1.305907972684991e+17, 1.305907972766244e+17, 1.305907972847496e+17, 1.30590797293031e+17, 1.305907973011562e+17, 1.305907973092814e+17, 1.305907973174067e+17, 1.305907973255319e+17, 1.305907973378758e+17, 1.305907973500639e+17, 1.305907973622516e+17, 1.305907973745957e+17, 1.305907973866272e+17, 1.305907973989713e+17, 1.305907974111592e+17, 1.305907974192844e+17, 1.305907974274097e+17, 1.305907974358473e+17, 1.305907974477226e+17, 1.305907974599104e+17, 1.305907974722546e+17, 1.305907974844424e+17, 1.305907974966303e+17, 1.30590797508818e+17, 1.305907975169432e+17, 1.305907975252247e+17, 1.305907975374125e+17, 1.305907975455377e+17, 1.305907975578817e+17, 1.305907975700695e+17, 1.305907975822574e+17, 1.305907975903827e+17, 1.305907976025705e+17, 1.305907976106957e+17, 1.30590797618821e+17, 1.305907976271023e+17, 1.305907976352276e+17, 1.305907976474154e+17, 1.305907976555406e+17, 1.305907976677285e+17, 1.305907976758537e+17, 1.305907976839789e+17, 1.305907976963229e+17, 1.305907977044483e+17, 1.305907977125734e+17, 1.305907977247612e+17, 1.305907977328864e+17, 1.305907977410117e+17, 1.305907977491369e+17, 1.305907977572621e+17, 1.305907977655436e+17, 1.305907977777315e+17, 1.305907977899192e+17, 1.30590797802107e+17, 1.305907978103885e+17, 1.305907978185137e+17, 1.305907978307016e+17, 1.30590797838983e+17, 1.305907978511708e+17, 1.305907978633587e+17, 1.305907978755465e+17, 1.305907978836717e+17, 1.30590797891797e+17, 1.305907979041411e+17, 1.30590797916329e+17, 1.305907979244541e+17, 1.305907979366419e+17, 1.305907979447671e+17, 1.305907979569549e+17, 1.305907979652364e+17, 1.305907979733617e+17, 1.305907979814868e+17, 1.30590797989612e+17, 1.305907979977372e+17, 1.305907980100814e+17, 1.305907980222692e+17, 1.305907980303944e+17, 1.305907980385197e+17, 1.305907980507075e+17, 1.305907980588326e+17, 1.305907980710205e+17, 1.30590798079302e+17, 1.305907980914898e+17, 1.305907981036776e+17, 1.305907981158655e+17, 1.305907981280532e+17, 1.305907981403973e+17, 1.305907981525851e+17, 1.30590798164773e+17, 1.305907981769608e+17, 1.305907981893048e+17, 1.305907982014926e+17, 1.305907982136805e+17, 1.305907982258684e+17, 1.305907982380562e+17, 1.30590798250244e+17, 1.305907982624317e+17, 1.305907982747758e+17, 1.305907982869637e+17, 1.305907982991515e+17, 1.305907983113394e+17, 1.305907983235272e+17, 1.305907983358712e+17, 1.305907983480591e+17, 1.305907983602469e+17, 1.305907983724348e+17, 1.305907983846226e+17, 1.305907983968104e+17, 1.305907984089983e+17, 1.305907984213423e+17, 1.305907984335302e+17, 1.305907984457179e+17, 1.305907984579058e+17, 1.305907984700937e+17, 1.305907984824376e+17, 1.305907984946255e+17, 1.305907985068133e+17, 1.305907985191574e+17, 1.305907985313453e+17, 1.305907985435331e+17, 1.305907985557208e+17, 1.305907985679086e+17, 1.305907985802528e+17, 1.305907985924406e+17, 1.305907986046285e+17, 1.305907986168163e+17, 1.30590798629004e+17, 1.305907986411919e+17, 1.305907986533797e+17, 1.305907986655675e+17, 1.305907986777554e+17, 1.305907986899432e+17, 1.305907987021311e+17, 1.305907987143188e+17, 1.305907987266629e+17, 1.305907987388508e+17, 1.305907987510385e+17, 1.305907987633827e+17, 1.305907987755704e+17, 1.305907987877583e+17, 1.305907988001024e+17, 1.305907988122902e+17, 1.30590798824478e+17, 1.305907988366659e+17, 1.305907988488538e+17, 1.305907988611977e+17, 1.305907988733856e+17, 1.305907988857295e+17, 1.305907988979176e+17, 1.305907989101053e+17, 1.305907989224494e+17, 1.305907989346372e+17, 1.30590798946825e+17, 1.30590798959169e+17, 1.305907989713569e+17, 1.305907989835448e+17, 1.305907989957325e+17, 1.305907990079204e+17, 1.305907990201083e+17, 1.305907990322961e+17, 1.30590799044484e+17, 1.305907990566717e+17, 1.305907990688595e+17, 1.305907990812036e+17, 1.305907990933914e+17, 1.305907991055793e+17, 1.30590799117767e+17, 1.305907991299549e+17, 1.30590799142299e+17, 1.305907991544868e+17, 1.30590799162612e+17, 1.305907991747999e+17, 1.305907991830813e+17, 1.305907991952691e+17, 1.30590799207457e+17, 1.305907992196448e+17, 1.305907992318326e+17, 1.305907992440205e+17, 1.305907992562083e+17, 1.305907992685523e+17, 1.305907992807402e+17, 1.30590799292928e+17, 1.305907993051159e+17, 1.3059079931746e+17, 1.305907993296477e+17, 1.305907993418355e+17, 1.305907993540234e+17, 1.305907993662112e+17, 1.305907993785553e+17, 1.305907993866806e+17, 1.305907993988684e+17, 1.305907994110561e+17, 1.30590799423244e+17, 1.305907994354318e+17, 1.305907994476196e+17, 1.305907994598075e+17, 1.305907994721516e+17, 1.305907994843395e+17, 1.305907994965272e+17, 1.30590799508715e+17, 1.305907995209029e+17, 1.305907995330907e+17, 1.305907995454348e+17, 1.305907995576225e+17, 1.305907995698104e+17, 1.305907995821544e+17, 1.305907995943423e+17, 1.3059079960653e+17, 1.305907996187178e+17, 1.30590799631062e+17, 1.305907996432498e+17, 1.305907996554377e+17, 1.305907996676255e+17, 1.305907996799697e+17, 1.305907996921573e+17, 1.305907997043452e+17, 1.305907997165331e+17, 1.305907997288771e+17, 1.30590799741065e+17, 1.30590799753409e+17, 1.305907997655968e+17, 1.305907997777847e+17, 1.305907997901288e+17, 1.305907998023165e+17, 1.305907998145044e+17, 1.305907998266922e+17, 1.305907998390363e+17, 1.305907998512242e+17, 1.30590799863412e+17, 1.305907998755999e+17, 1.305907998879438e+17, 1.305907999001317e+17, 1.305907999123195e+17, 1.305907999245073e+17, 1.305907999366952e+17, 1.305907999488829e+17, 1.30590799961227e+17, 1.305907999734149e+17, 1.305907999856027e+17, 1.305907999977905e+17, 1.305908000099782e+17, 1.305908000223224e+17, 1.305908000345102e+17, 1.305908000466981e+17, 1.305908000588859e+17, 1.305908000710737e+17, 1.305908000834179e+17, 1.305908000956056e+17, 1.305908001077935e+17, 1.305908001199813e+17, 1.305908001323254e+17, 1.305908001445133e+17, 1.305908001567011e+17, 1.305908001688888e+17, 1.305908001812329e+17, 1.305908001934207e+17, 1.305908002056086e+17, 1.305908002177964e+17, 1.305908002301404e+17, 1.305908002423283e+17, 1.305908002545161e+17, 1.305908002667039e+17, 1.305908002788918e+17, 1.305908002912358e+17, 1.305908003034237e+17, 1.305908003156115e+17, 1.305908003279556e+17, 1.305908003401435e+17, 1.305908003523313e+17, 1.30590800364519e+17, 1.30590800376863e+17, 1.30590800389051e+17, 1.305908004012388e+17, 1.305908004134266e+17, 1.305908004256145e+17, 1.305908004378022e+17, 1.3059080044999e+17, 1.305908004623341e+17, 1.30590800474522e+17, 1.305908004867098e+17, 1.305908004988975e+17, 1.305908005110854e+17, 1.305908005234295e+17, 1.305908005356174e+17, 1.305908005478052e+17, 1.30590800559993e+17, 1.305908005721809e+17, 1.305908005843686e+17, 1.305908005967128e+17, 1.305908006089006e+17, 1.305908006210884e+17, 1.305908006332762e+17, 1.305908006454641e+17, 1.305908006576518e+17, 1.305908006698397e+17, 1.305908006821838e+17, 1.305908006943715e+17, 1.305908007065594e+17, 1.305908007187473e+17, 1.30590800730935e+17, 1.305908007431228e+17, 1.305908007554669e+17, 1.305908007676548e+17, 1.305908007798427e+17, 1.305908007920303e+17, 1.305908008042182e+17, 1.305908008165623e+17, 1.305908008287501e+17, 1.30590800840938e+17, 1.305908008531258e+17, 1.3059080086547e+17, 1.305908008776577e+17, 1.305908008898455e+17, 1.305908009020334e+17, 1.305908009143775e+17, 1.305908009265652e+17, 1.30590800938753e+17, 1.305908009509409e+17, 1.305908009631287e+17, 1.305908009754728e+17, 1.305908009876605e+17, 1.305908009998484e+17, 1.305908010120364e+17, 1.305908010242241e+17, 1.305908010364119e+17, 1.305908010485997e+17, 1.305908010609439e+17, 1.305908010731316e+17, 1.305908010853194e+17, 1.305908010975073e+17, 1.305908011096951e+17, 1.305908011220393e+17, 1.305908011342271e+17, 1.305908011464148e+17, 1.305908011586028e+17, 1.305908011707905e+17, 1.305908011829783e+17, 1.305908011951662e+17, 1.305908012075103e+17, 1.30590801219698e+17, 1.305908012320421e+17, 1.3059080124423e+17, 1.305908012564177e+17, 1.305908012686056e+17, 1.305908012807935e+17, 1.305908012931375e+17, 1.305908013053253e+17, 1.305908013175131e+17, 1.30590801329701e+17, 1.305908013418888e+17, 1.305908013540765e+17, 1.305908013664207e+17, 1.305908013786085e+17, 1.305908013907964e+17, 1.305908014029842e+17, 1.30590801415172e+17, 1.30590801427516e+17, 1.305908014397039e+17, 1.305908014518918e+17, 1.305908014640796e+17, 1.305908014762674e+17, 1.305908014884552e+17, 1.305908015006429e+17, 1.305908015129871e+17, 1.305908015251749e+17, 1.305908015373628e+17, 1.305908015497068e+17, 1.305908015618947e+17, 1.305908015740824e+17, 1.305908015862703e+17, 1.305908015986144e+17, 1.305908016108022e+17, 1.305908016229901e+17, 1.305908016351779e+17, 1.30590801647522e+17, 1.305908016597098e+17, 1.305908016718976e+17, 1.305908016840854e+17, 1.305908016962732e+17, 1.305908017086173e+17, 1.305908017208051e+17, 1.30590801732993e+17, 1.305908017451808e+17, 1.305908017573686e+17, 1.305908017695565e+17, 1.305908017817443e+17, 1.305908017940883e+17, 1.305908018062761e+17, 1.30590801818464e+17, 1.305908018308081e+17, 1.305908018429958e+17, 1.305908018551837e+17, 1.305908018673715e+17, 1.305908018797157e+17, 1.305908018919035e+17, 1.305908019040913e+17, 1.305908019162792e+17, 1.305908019284669e+17, 1.30590801940811e+17, 1.305908019529988e+17, 1.305908019651867e+17, 1.305908019773745e+17, 1.305908019895622e+17, 1.305908020017501e+17, 1.305908020139379e+17, 1.305908020262821e+17, 1.305908020384698e+17, 1.305908020506577e+17, 1.305908020628454e+17, 1.305908020751896e+17, 1.305908020873774e+17, 1.305908020995652e+17, 1.305908021117531e+17, 1.305908021239409e+17, 1.305908021362851e+17, 1.305908021484728e+17, 1.305908021606606e+17, 1.305908021728485e+17, 1.305908021851924e+17, 1.305908021973805e+17, 1.30590802209412e+17, 1.305908022217559e+17, 1.305908022339438e+17, 1.305908022461316e+17, 1.305908022583195e+17, 1.305908022706636e+17, 1.305908022826952e+17, 1.305908022950392e+17, 1.30590802307227e+17, 1.305908023194149e+17, 1.305908023317588e+17, 1.305908023439468e+17, 1.305908023561345e+17, 1.305908023683223e+17, 1.305908023805102e+17, 1.305908023928543e+17, 1.305908024050422e+17, 1.3059080241723e+17, 1.305908024294177e+17, 1.305908024416056e+17, 1.305908024537934e+17, 1.305908024661376e+17, 1.305908024783252e+17, 1.305908024905132e+17, 1.305908025027011e+17, 1.305908025148888e+17, 1.305908025270767e+17, 1.305908025394207e+17, 1.305908025516086e+17, 1.305908025637964e+17, 1.305908025759841e+17, 1.30590802588172e+17, 1.30590802600516e+17, 1.305908026127039e+17, 1.305908026248916e+17, 1.305908026370796e+17, 1.305908026494236e+17, 1.305908026616114e+17, 1.305908026739555e+17, 1.305908026861434e+17, 1.305908026983313e+17, 1.30590802710519e+17, 1.305908027227068e+17, 1.305908027348947e+17, 1.305908027472388e+17, 1.305908027594266e+17, 1.305908027716143e+17, 1.305908027838022e+17, 1.305908027961462e+17, 1.305908028083341e+17, 1.30590802820522e+17, 1.305908028327098e+17, 1.305908028448975e+17, 1.305908028570853e+17, 1.305908028692732e+17, 1.305908028814611e+17, 1.305908028938052e+17, 1.30590802905993e+17, 1.305908029181807e+17, 1.305908029303686e+17, 1.305908029425564e+17, 1.305908029547442e+17, 1.305908029670884e+17, 1.305908029792762e+17, 1.305908029914641e+17, 1.30590803003808e+17, 1.305908030159959e+17, 1.305908030281837e+17, 1.305908030405277e+17, 1.305908030527155e+17, 1.305908030649034e+17, 1.305908030770913e+17, 1.305908030892791e+17, 1.305908031016232e+17, 1.305908031138109e+17, 1.305908031259988e+17, 1.305908031383429e+17, 1.305908031505307e+17, 1.305908031627186e+17, 1.305908031749064e+17, 1.305908031872506e+17, 1.305908031994383e+17, 1.305908032116261e+17, 1.305908032238139e+17, 1.305908032360017e+17, 1.305908032481896e+17, 1.305908032603775e+17, 1.305908032727215e+17, 1.305908032849093e+17, 1.305908032970971e+17, 1.30590803309285e+17, 1.305908033214728e+17, 1.305908033336607e+17, 1.305908033460046e+17, 1.305908033581925e+17, 1.305908033703803e+17, 1.305908033825681e+17, 1.30590803394756e+17, 1.305908034069437e+17, 1.305908034191316e+17, 1.305908034313194e+17, 1.305908034435072e+17, 1.305908034556951e+17, 1.305908034678829e+17, 1.305908034800707e+17, 1.305908034922586e+17, 1.305908035046026e+17, 1.305908035167905e+17, 1.305908035289783e+17, 1.305908035413224e+17, 1.30590803553354e+17, 1.305908035655418e+17, 1.30590803577886e+17, 1.305908035900737e+17, 1.305908036022615e+17, 1.305908036146056e+17, 1.305908036267935e+17, 1.305908036389812e+17, 1.30590803651169e+17, 1.305908036635131e+17, 1.305908036757009e+17, 1.305908036878888e+17, 1.305908037000767e+17, 1.305908037122643e+17, 1.305908037244522e+17, 1.3059080373664e+17, 1.305908037489842e+17, 1.30590803761172e+17, 1.305908037733597e+17, 1.305908037855476e+17, 1.305908037977354e+17, 1.305908038099233e+17, 1.305908038222674e+17, 1.305908038344552e+17, 1.305908038466431e+17, 1.305908038588308e+17, 1.305908038710188e+17, 1.305908038833627e+17, 1.305908038955506e+17, 1.305908039077384e+17, 1.305908039199261e+17, 1.305908039322703e+17, 1.305908039444581e+17, 1.30590803956646e+17, 1.305908039688337e+17, 1.305908039811779e+17, 1.305908039933656e+17, 1.305908040055534e+17, 1.305908040177413e+17, 1.305908040300854e+17, 1.305908040422733e+17, 1.305908040544611e+17, 1.305908040666488e+17, 1.305908040788367e+17, 1.305908040911808e+17, 1.305908041033686e+17, 1.305908041155565e+17, 1.305908041277443e+17, 1.305908041399322e+17, 1.305908041522762e+17, 1.30590804164464e+17, 1.305908041766518e+17, 1.305908041889958e+17, 1.305908042011836e+17, 1.305908042133715e+17, 1.305908042255593e+17, 1.305908042377472e+17, 1.305908042500913e+17, 1.30590804262279e+17, 1.305908042744669e+17, 1.305908042866547e+17, 1.305908042988426e+17, 1.305908043110304e+17, 1.305908043232182e+17, 1.305908043354061e+17, 1.3059080434775e+17, 1.30590804359938e+17, 1.305908043721258e+17, 1.305908043843136e+17, 1.305908043965015e+17, 1.305908044088454e+17, 1.305908044210333e+17, 1.305908044332211e+17, 1.305908044454089e+17, 1.30590804457753e+17, 1.305908044699409e+17, 1.305908044821286e+17, 1.305908044944727e+17, 1.305908045065043e+17, 1.305908045188484e+17, 1.305908045310363e+17, 1.305908045432241e+17, 1.305908045554118e+17, 1.305908045675997e+17, 1.305908045797875e+17, 1.305908045919753e+17, 1.305908046043194e+17, 1.305908046165073e+17, 1.305908046286952e+17, 1.305908046410391e+17, 1.30590804653227e+17, 1.305908046654148e+17, 1.305908046776027e+17, 1.305908046897905e+17, 1.305908047021345e+17, 1.305908047143224e+17, 1.305908047265101e+17, 1.305908047386981e+17, 1.305908047508859e+17, 1.3059080476323e+17, 1.305908047754177e+17, 1.305908047876055e+17, 1.305908047997934e+17, 1.305908048119812e+17, 1.305908048243254e+17, 1.305908048365132e+17, 1.305908048487009e+17, 1.305908048610451e+17, 1.305908048732328e+17, 1.305908048854207e+17, 1.305908048976084e+17, 1.305908049097964e+17, 1.305908049221404e+17, 1.305908049343282e+17, 1.305908049465161e+17, 1.305908049587039e+17, 1.305908049708916e+17, 1.305908049830796e+17, 1.305908049954236e+17, 1.305908050076114e+17, 1.305908050197992e+17, 1.305908050319871e+17, 1.305908050441748e+17, 1.305908050563628e+17, 1.305908050687068e+17, 1.305908050808946e+17, 1.305908050930825e+17, 1.305908051052703e+17, 1.305908051174582e+17, 1.305908051298022e+17, 1.3059080514199e+17, 1.305908051541778e+17, 1.305908051663657e+17, 1.305908051785536e+17, 1.305908051908975e+17, 1.305908052030854e+17, 1.305908052152732e+17, 1.305908052276174e+17, 1.305908052398052e+17, 1.30590805251993e+17, 1.305908052641807e+17, 1.305908052763685e+17, 1.305908052887127e+17, 1.305908053009005e+17, 1.305908053130884e+17, 1.305908053252762e+17, 1.305908053374639e+17, 1.305908053496518e+17, 1.305908053618396e+17, 1.305908053741838e+17, 1.305908053863716e+17, 1.305908053985592e+17, 1.305908054107473e+17, 1.30590805422935e+17, 1.305908054352791e+17, 1.305908054474669e+17, 1.305908054596547e+17, 1.305908054718426e+17, 1.305908054840303e+17, 1.305908054962182e+17, 1.305908055085623e+17, 1.305908055207501e+17, 1.30590805532938e+17, 1.305908055451258e+17, 1.305908055573137e+17, 1.305908055695014e+17, 1.305908055818455e+17, 1.305908055940333e+17, 1.305908056062211e+17, 1.30590805618409e+17, 1.30590805630753e+17, 1.305908056429409e+17, 1.305908056551287e+17, 1.305908056673165e+17, 1.305908056796605e+17, 1.305908056918484e+17, 1.305908057040362e+17, 1.30590805716224e+17, 1.305908057284119e+17, 1.30590805740756e+17, 1.305908057529439e+17, 1.305908057651316e+17, 1.305908057773194e+17, 1.305908057895073e+17, 1.305908058018513e+17, 1.305908058140392e+17, 1.305908058262269e+17, 1.305908058384147e+17, 1.305908058506026e+17, 1.305908058627904e+17, 1.305908058751346e+17, 1.305908058873224e+17, 1.305908058995101e+17, 1.30590805911698e+17, 1.305908059238858e+17, 1.305908059360737e+17, 1.305908059484177e+17, 1.305908059606056e+17, 1.305908059727935e+17, 1.305908059849812e+17, 1.30590805997169e+17, 1.305908060095131e+17, 1.30590806021701e+17, 1.305908060338888e+17, 1.30590806046233e+17, 1.305908060584206e+17, 1.305908060706085e+17, 1.305908060827963e+17, 1.305908060949842e+17, 1.30590806107172e+17, 1.30590806119516e+17, 1.305908061317039e+17, 1.305908061438917e+17, 1.305908061560795e+17, 1.305908061682674e+17, 1.305908061804552e+17, 1.305908061926429e+17, 1.30590806204987e+17, 1.305908062171749e+17, 1.305908062293628e+17, 1.305908062415506e+17, 1.305908062537384e+17, 1.305908062660824e+17, 1.305908062782702e+17, 1.305908062904581e+17, 1.305908063026459e+17, 1.305908063148338e+17, 1.305908063271777e+17, 1.305908063393656e+17, 1.305908063515535e+17, 1.305908063637412e+17, 1.305908063759291e+17, 1.305908063881169e+17, 1.305908064004611e+17, 1.305908064126488e+17, 1.305908064248366e+17, 1.305908064371808e+17, 1.305908064492123e+17, 1.305908064615565e+17, 1.305908064737443e+17, 1.30590806485932e+17, 1.305908064981199e+17, 1.305908065103077e+17, 1.305908065224956e+17, 1.305908065346834e+17, 1.305908065470275e+17, 1.305908065592152e+17, 1.30590806571403e+17, 1.305908065837472e+17, 1.30590806595935e+17, 1.305908066081229e+17, 1.305908066203107e+17, 1.305908066324984e+17, 1.305908066448425e+17, 1.305908066570304e+17, 1.305908066692182e+17, 1.30590806681406e+17, 1.305908066935939e+17, 1.305908067057816e+17, 1.305908067181258e+17, 1.305908067303136e+17, 1.305908067425014e+17, 1.305908067546893e+17, 1.305908067668771e+17, 1.305908067792212e+17, 1.30590806791409e+17, 1.305908068035967e+17, 1.305908068157846e+17, 1.305908068281286e+17, 1.305908068403165e+17, 1.305908068525043e+17, 1.305908068646921e+17, 1.3059080687688e+17, 1.305908068892241e+17, 1.30590806901412e+17, 1.305908069135997e+17, 1.305908069257875e+17, 1.305908069379753e+17, 1.305908069503195e+17, 1.305908069625073e+17, 1.30590806974695e+17, 1.305908069868829e+17, 1.30590806999227e+17, 1.305908070114149e+17, 1.305908070236027e+17, 1.305908070357905e+17, 1.305908070479784e+17, 1.305908070601661e+17, 1.305908070723539e+17, 1.30590807084698e+17, 1.305908070968859e+17, 1.305908071090737e+17, 1.305908071212614e+17, 1.305908071334493e+17, 1.305908071456371e+17, 1.305908071578249e+17, 1.305908071701691e+17, 1.305908071823567e+17, 1.305908071945446e+17, 1.305908072067325e+17, 1.305908072189203e+17, 1.305908072311081e+17, 1.305908072434522e+17, 1.305908072556401e+17, 1.305908072678278e+17, 1.305908072800157e+17, 1.305908072922035e+17, 1.305908073045476e+17, 1.305908073167355e+17, 1.305908073290796e+17, 1.305908073411112e+17, 1.305908073532989e+17, 1.30590807365643e+17, 1.305908073778308e+17, 1.305908073900187e+17, 1.305908074022066e+17, 1.305908074143944e+17, 1.305908074265821e+17, 1.305908074389262e+17, 1.30590807451114e+17, 1.305908074633019e+17, 1.305908074754897e+17, 1.305908074876776e+17, 1.305908074998653e+17, 1.305908075122094e+17, 1.305908075243972e+17, 1.30590807536585e+17, 1.305908075489292e+17, 1.305908075611169e+17, 1.305908075733048e+17, 1.305908075854926e+17, 1.305908075976804e+17, 1.305908076100244e+17, 1.305908076222122e+17, 1.305908076344003e+17, 1.30590807646588e+17, 1.305908076587758e+17, 1.305908076709636e+17, 1.305908076833076e+17, 1.305908076954956e+17, 1.305908077076833e+17, 1.305908077198712e+17, 1.305908077322152e+17, 1.305908077444031e+17, 1.30590807756591e+17, 1.305908077687786e+17, 1.305908077809665e+17, 1.305908077933106e+17, 1.305908078053422e+17, 1.305908078176863e+17, 1.30590807829874e+17, 1.30590807842062e+17, 1.30590807854406e+17, 1.305908078665938e+17, 1.305908078787817e+17, 1.305908078909695e+17, 1.305908079031574e+17, 1.305908079153452e+17, 1.305908079275331e+17, 1.305908079397208e+17, 1.305908079519086e+17, 1.305908079640965e+17, 1.305908079762843e+17, 1.305908079886284e+17, 1.305908080008161e+17, 1.30590808013004e+17, 1.305908080251918e+17, 1.305908080373796e+17, 1.305908080495675e+17, 1.305908080619116e+17, 1.305908080740995e+17, 1.305908080862872e+17, 1.305908080984749e+17, 1.305908081106628e+17, 1.305908081228507e+17, 1.305908081350385e+17, 1.305908081472264e+17, 1.305908081594141e+17, 1.305908081717582e+17, 1.30590808183946e+17, 1.305908081961339e+17, 1.305908082083217e+17, 1.305908082205094e+17, 1.305908082326973e+17, 1.305908082450414e+17, 1.305908082572293e+17, 1.305908082694171e+17, 1.305908082816049e+17, 1.305908082937928e+17, 1.305908083059805e+17, 1.305908083181683e+17, 1.305908083305124e+17, 1.305908083427003e+17, 1.305908083548881e+17, 1.305908083670758e+17, 1.3059080837942e+17, 1.305908083916077e+17, 1.305908084037957e+17, 1.305908084159835e+17, 1.305908084281713e+17, 1.305908084403592e+17, 1.305908084525468e+17, 1.30590808464891e+17, 1.305908084770788e+17, 1.305908084892667e+17, 1.305908085014545e+17, 1.305908085136422e+17, 1.305908085258301e+17, 1.305908085381742e+17, 1.305908085503621e+17, 1.305908085625499e+17, 1.305908085747377e+17, 1.305908085869256e+17, 1.305908085991133e+17, 1.305908086114574e+17, 1.305908086236452e+17, 1.305908086359892e+17, 1.30590808648177e+17, 1.305908086602086e+17, 1.305908086723965e+17, 1.305908086847406e+17, 1.305908086969284e+17, 1.305908087091162e+17, 1.305908087213039e+17, 1.305908087334918e+17, 1.305908087456797e+17, 1.305908087578675e+17, 1.305908087702116e+17, 1.305908087823994e+17, 1.305908087945873e+17, 1.30590808806775e+17, 1.305908088189629e+17, 1.30590808831307e+17, 1.305908088434948e+17, 1.305908088556826e+17, 1.305908088680268e+17, 1.305908088802145e+17, 1.305908088922461e+17, 1.305908089044339e+17, 1.30590808916778e+17, 1.305908089289658e+17, 1.305908089413098e+17, 1.305908089534977e+17, 1.305908089656855e+17, 1.305908089778733e+17, 1.305908089900612e+17, 1.305908090024052e+17, 1.30590809014593e+17, 1.305908090267809e+17, 1.305908090389687e+17, 1.305908090511566e+17, 1.305908090635005e+17, 1.305908090756884e+17, 1.305908090878764e+17, 1.305908091002204e+17, 1.305908091122519e+17, 1.305908091244397e+17, 1.305908091367839e+17, 1.305908091489716e+17, 1.305908091611594e+17, 1.305908091733473e+17, 1.305908091856914e+17, 1.305908091978792e+17, 1.305908092100669e+17, 1.305908092222548e+17, 1.305908092345989e+17, 1.305908092467868e+17, 1.305908092589746e+17, 1.305908092711624e+17, 1.305908092833503e+17, 1.305908092956943e+17, 1.305908093078822e+17, 1.305908093200699e+17, 1.305908093322578e+17, 1.305908093444456e+17, 1.305908093566335e+17, 1.305908093689775e+17, 1.305908093811653e+17, 1.305908093933532e+17, 1.30590809405541e+17, 1.305908094177288e+17, 1.305908094299167e+17, 1.305908094422606e+17, 1.305908094544485e+17, 1.305908094666363e+17, 1.305908094788241e+17, 1.30590809491012e+17, 1.30590809503356e+17, 1.305908095155439e+17, 1.305908095277317e+17, 1.305908095399195e+17, 1.305908095521074e+17, 1.305908095642952e+17, 1.305908095764831e+17, 1.30590809588827e+17, 1.305908096010149e+17, 1.305908096132027e+17, 1.305908096253906e+17, 1.305908096375785e+17, 1.305908096497661e+17, 1.305908096621102e+17, 1.30590809674298e+17, 1.305908096864859e+17, 1.305908096986738e+17, 1.305908097108616e+17, 1.305908097232056e+17, 1.305908097353934e+17, 1.305908097475813e+17, 1.305908097599254e+17, 1.305908097721133e+17, 1.305908097843011e+17, 1.305908097964888e+17, 1.305908098086767e+17, 1.305908098210207e+17, 1.305908098332086e+17, 1.305908098453965e+17, 1.305908098575841e+17, 1.30590809869772e+17, 1.305908098819598e+17, 1.30590809894304e+17, 1.305908099064918e+17, 1.305908099186796e+17, 1.305908099308673e+17, 1.305908099430551e+17, 1.30590809955243e+17, 1.305908099675871e+17, 1.30590809979775e+17, 1.305908099919628e+17, 1.305908100041505e+17, 1.305908100163384e+17, 1.305908100286825e+17, 1.305908100408704e+17, 1.305908100530582e+17, 1.305908100654022e+17, 1.3059081007759e+17, 1.305908100897779e+17, 1.305908101019657e+17, 1.305908101143098e+17, 1.305908101264975e+17, 1.305908101386853e+17, 1.305908101508732e+17, 1.305908101630611e+17, 1.305908101754052e+17, 1.30590810187593e+17, 1.305908101997807e+17, 1.305908102119686e+17, 1.305908102241564e+17, 1.305908102365006e+17, 1.305908102486884e+17, 1.305908102610324e+17, 1.305908102732202e+17, 1.30590810285408e+17, 1.305908102975959e+17, 1.305908103097837e+17, 1.305908103221279e+17, 1.305908103343156e+17, 1.305908103465034e+17, 1.305908103586912e+17, 1.30590810370879e+17, 1.30590810383067e+17, 1.305908103954109e+17, 1.305908104075988e+17, 1.305908104199428e+17, 1.305908104321307e+17, 1.305908104443186e+17, 1.305908104565064e+17, 1.305908104688504e+17, 1.305908104810382e+17, 1.305908104932261e+17, 1.305908105054139e+17, 1.305908105177581e+17, 1.305908105299457e+17, 1.305908105421336e+17, 1.305908105543214e+17, 1.305908105665092e+17, 1.305908105788534e+17, 1.305908105910412e+17, 1.305908106032291e+17, 1.30590810615573e+17, 1.305908106277609e+17, 1.305908106399487e+17, 1.305908106521366e+17, 1.305908106643245e+17, 1.305908106726058e+17, 1.305908106847936e+17, 1.305908106969815e+17, 1.305908107091693e+17, 1.305908107213571e+17, 1.305908107337012e+17, 1.30590810745889e+17, 1.305908107540142e+17, 1.305908107662021e+17, 1.305908107783899e+17, 1.305908107905777e+17, 1.305908108029217e+17, 1.305908108151096e+17, 1.305908108272974e+17, 1.305908108396415e+17, 1.305908108518294e+17, 1.305908108640172e+17, 1.305908108762051e+17, 1.30590810888549e+17, 1.305908109007369e+17, 1.305908109088621e+17, 1.3059081092105e+17, 1.30590810933394e+17, 1.305908109455818e+17, 1.305908109537071e+17, 1.305908109660511e+17, 1.30590810978239e+17, 1.305908109904269e+17, 1.305908110026145e+17, 1.305908110148024e+17, 1.305908110271465e+17, 1.305908110393343e+17, 1.30590811051522e+17, 1.3059081106371e+17, 1.305908110758977e+17, 1.305908110882419e+17, 1.305908111004297e+17, 1.305908111126175e+17, 1.305908111249617e+17, 1.305908111371494e+17, 1.305908111493373e+17, 1.305908111615251e+17, 1.305908111738692e+17, 1.30590811186057e+17, 1.305908111982447e+17, 1.305908112104326e+17, 1.305908112226204e+17, 1.305908112348083e+17, 1.305908112471523e+17, 1.305908112593402e+17, 1.305908112715279e+17, 1.305908112837157e+17, 1.305908112959036e+17, 1.305908113080914e+17, 1.305908113204356e+17, 1.305908113326234e+17, 1.305908113448111e+17, 1.30590811356999e+17, 1.305908113691868e+17, 1.305908113813747e+17, 1.305908113935625e+17, 1.305908114059066e+17, 1.305908114180945e+17, 1.305908114302821e+17, 1.305908114423137e+17, 1.305908114546579e+17, 1.305908114668457e+17, 1.305908114790336e+17, 1.305908114913775e+17, 1.305908115035654e+17, 1.305908115155969e+17, 1.30590811527941e+17, 1.305908115401289e+17, 1.305908115523167e+17, 1.305908115646607e+17, 1.305908115768485e+17, 1.305908115890364e+17, 1.305908116012242e+17, 1.30590811613412e+17, 1.305908116255999e+17, 1.305908116377876e+17, 1.305908116501318e+17, 1.305908116623196e+17, 1.305908116745074e+17, 1.305908116866953e+17, 1.305908116990394e+17, 1.305908117112271e+17, 1.30590811723415e+17, 1.305908117356028e+17, 1.305908117477907e+17, 1.305908117599784e+17, 1.305908117723226e+17, 1.305908117845103e+17, 1.305908117966982e+17, 1.30590811808886e+17, 1.305908118210738e+17, 1.305908118332616e+17, 1.305908118456056e+17, 1.305908118577935e+17, 1.305908118699813e+17, 1.305908118823255e+17, 1.305908118945133e+17, 1.305908119067011e+17, 1.30590811918889e+17, 1.30590811931233e+17, 1.305908119434208e+17, 1.305908119556086e+17, 1.305908119677965e+17, 1.305908119799843e+17, 1.305908119923284e+17, 1.305908120045162e+17, 1.30590812016704e+17, 1.305908120288919e+17, 1.305908120410797e+17, 1.305908120532675e+17, 1.305908120656115e+17, 1.305908120777994e+17, 1.305908120899872e+17, 1.30590812102175e+17, 1.305908121143629e+17, 1.305908121267069e+17, 1.305908121388948e+17, 1.305908121510826e+17, 1.305908121632704e+17, 1.305908121754583e+17, 1.305908121876461e+17, 1.305908121998339e+17, 1.305908122121779e+17, 1.305908122243657e+17, 1.305908122365536e+17, 1.305908122487414e+17, 1.305908122609293e+17, 1.305908122731172e+17, 1.305908122854611e+17, 1.30590812297649e+17, 1.305908123098367e+17, 1.305908123220246e+17, 1.305908123343686e+17, 1.305908123465565e+17, 1.305908123587443e+17, 1.305908123710885e+17, 1.305908123832762e+17, 1.305908123954641e+17, 1.30590812407652e+17, 1.305908124198397e+17, 1.305908124320275e+17, 1.305908124443716e+17, 1.305908124565595e+17, 1.305908124687473e+17, 1.30590812480935e+17, 1.305908124931229e+17, 1.305908125053107e+17, 1.305908125176548e+17, 1.305908125298426e+17, 1.305908125420305e+17, 1.305908125542184e+17, 1.305908125664061e+17, 1.305908125787502e+17, 1.30590812590938e+17, 1.305908126031259e+17, 1.305908126153137e+17, 1.305908126276577e+17, 1.305908126398456e+17, 1.305908126520334e+17, 1.305908126642213e+17, 1.305908126764091e+17, 1.305908126887532e+17, 1.305908127009409e+17, 1.305908127131287e+17, 1.305908127253166e+17, 1.305908127376605e+17, 1.305908127498486e+17, 1.305908127620364e+17, 1.305908127742241e+17, 1.305908127864119e+17, 1.30590812798756e+17, 1.305908128109439e+17, 1.305908128231316e+17, 1.305908128353196e+17, 1.305908128475073e+17, 1.305908128596951e+17, 1.30590812871883e+17, 1.305908128842271e+17, 1.30590812896415e+17, 1.305908129086028e+17, 1.305908129207905e+17, 1.305908129329783e+17, 1.305908129453224e+17, 1.305908129575103e+17, 1.30590812969698e+17, 1.305908129820421e+17, 1.305908129942299e+17, 1.305908130064178e+17, 1.305908130186057e+17, 1.305908130307933e+17, 1.305908130431375e+17, 1.305908130553253e+17, 1.305908130675132e+17, 1.30590813079701e+17, 1.305908130918888e+17, 1.305908131040767e+17, 1.305908131164207e+17, 1.305908131286085e+17, 1.305908131407964e+17, 1.305908131529842e+17, 1.305908131651721e+17, 1.305908131773599e+17, 1.305908131897039e+17, 1.305908132018917e+17, 1.305908132140796e+17, 1.305908132262674e+17, 1.305908132384552e+17, 1.305908132506431e+17, 1.30590813262987e+17, 1.305908132751749e+17, 1.305908132873627e+17, 1.305908132995506e+17, 1.305908133117384e+17, 1.305908133239261e+17, 1.305908133362703e+17, 1.305908133484581e+17, 1.30590813360646e+17, 1.305908133728338e+17, 1.305908133850216e+17, 1.305908133973656e+17, 1.305908134095534e+17, 1.305908134217414e+17, 1.305908134339292e+17, 1.30590813446117e+17, 1.305908134583048e+17, 1.305908134704925e+17, 1.305908134828367e+17, 1.305908134950245e+17, 1.305908135073686e+17, 1.305908135195564e+17, 1.305908135317443e+17, 1.30590813543932e+17, 1.305908135561198e+17, 1.30590813568464e+17, 1.305908135806518e+17, 1.305908135928397e+17, 1.305908136050275e+17, 1.305908136173715e+17, 1.305908136295594e+17, 1.305908136417472e+17, 1.30590813653935e+17, 1.305908136661228e+17, 1.305908136784669e+17, 1.305908136906547e+17, 1.305908137028425e+17, 1.305908137150304e+17, 1.305908137273745e+17, 1.305908137395622e+17, 1.3059081375175e+17, 1.305908137639379e+17, 1.305908137761257e+17, 1.305908137883135e+17, 1.305908138006577e+17, 1.305908138128454e+17, 1.305908138250333e+17, 1.305908138372211e+17, 1.305908138494089e+17, 1.30590813861753e+17, 1.305908138737846e+17, 1.305908138861288e+17, 1.305908138983164e+17, 1.305908139105043e+17, 1.305908139226921e+17, 1.305908139350362e+17, 1.305908139472239e+17, 1.305908139594118e+17, 1.305908139715997e+17, 1.305908139837874e+17, 1.305908139959753e+17, 1.305908140081632e+17, 1.305908140205071e+17, 1.30590814032695e+17, 1.305908140448828e+17, 1.305908140570707e+17, 1.305908140692585e+17, 1.305908140814463e+17, 1.305908140936342e+17, 1.30590814105822e+17, 1.305908141180097e+17, 1.305908141301976e+17, 1.305908141425417e+17, 1.305908141547296e+17, 1.305908141669174e+17, 1.305908141792614e+17, 1.305908141912931e+17, 1.305908142034808e+17, 1.305908142156687e+17, 1.305908142280128e+17, 1.305908142402006e+17, 1.305908142525446e+17, 1.305908142647324e+17, 1.305908142769202e+17, 1.30590814289108e+17, 1.30590814301296e+17, 1.305908143134838e+17, 1.305908143258278e+17, 1.305908143378593e+17, 1.305908143500471e+17, 1.305908143623913e+17, 1.305908143745791e+17, 1.30590814386767e+17, 1.30590814399111e+17, 1.305908144112988e+17, 1.305908144234867e+17, 1.305908144356745e+17, 1.305908144480186e+17, 1.305908144602063e+17, 1.305908144725504e+17, 1.305908144847382e+17, 1.305908144969262e+17, 1.30590814509114e+17, 1.305908145213018e+17, 1.305908145334895e+17, 1.305908145456773e+17, 1.305908145580215e+17, 1.305908145702093e+17, 1.305908145823972e+17, 1.30590814594585e+17, 1.30590814606929e+17, 1.305908146191169e+17, 1.305908146313047e+17, 1.305908146434926e+17, 1.305908146556804e+17, 1.305908146680244e+17, 1.305908146802122e+17, 1.305908146924e+17, 1.305908147045879e+17, 1.305908147167757e+17, 1.305908147289636e+17, 1.305908147413075e+17, 1.305908147534954e+17, 1.305908147656833e+17, 1.305908147778711e+17, 1.305908147900589e+17, 1.305908148024029e+17, 1.305908148145908e+17, 1.305908148267786e+17, 1.305908148389664e+17, 1.305908148513106e+17, 1.305908148634984e+17, 1.305908148756863e+17, 1.30590814887874e+17, 1.305908149002181e+17, 1.305908149124059e+17, 1.305908149245937e+17, 1.305908149367816e+17, 1.305908149489693e+17, 1.305908149611572e+17, 1.305908149735012e+17, 1.305908149856891e+17, 1.305908149978769e+17, 1.305908150100646e+17, 1.305908150222525e+17, 1.305908150345966e+17, 1.305908150467845e+17, 1.305908150589723e+17, 1.305908150713164e+17, 1.305908150835041e+17, 1.30590815095692e+17, 1.305908151078799e+17, 1.305908151202239e+17, 1.305908151324118e+17, 1.305908151445996e+17, 1.305908151567873e+17, 1.305908151689752e+17, 1.305908151813193e+17, 1.305908151935071e+17, 1.305908152056948e+17, 1.30590815218039e+17, 1.305908152302268e+17, 1.305908152424147e+17, 1.305908152547588e+17, 1.305908152669466e+17, 1.305908152791343e+17, 1.305908152913221e+17, 1.305908153035101e+17, 1.305908153156979e+17, 1.305908153278857e+17, 1.305908153402298e+17, 1.305908153524175e+17, 1.305908153646054e+17, 1.305908153767932e+17, 1.305908153889811e+17, 1.305908154011689e+17, 1.30590815413513e+17, 1.305908154257007e+17, 1.305908154378885e+17, 1.305908154500764e+17, 1.305908154622642e+17, 1.305908154746084e+17, 1.305908154867962e+17, 1.305908154989839e+17, 1.305908155111718e+17, 1.305908155233596e+17, 1.305908155355475e+17, 1.305908155478915e+17, 1.305908155600794e+17, 1.305908155722673e+17, 1.30590815584455e+17, 1.305908155966428e+17, 1.305908156088306e+17, 1.305908156211747e+17, 1.305908156333626e+17, 1.305908156455503e+17, 1.305908156577382e+17, 1.30590815669926e+17, 1.305908156821138e+17, 1.305908156944579e+17, 1.305908157066458e+17, 1.305908157188335e+17, 1.305908157310213e+17, 1.305908157432092e+17, 1.305908157555533e+17, 1.305908157677412e+17, 1.30590815779929e+17, 1.305908157921167e+17, 1.305908158044608e+17, 1.305908158166486e+17, 1.305908158288365e+17, 1.305908158410244e+17, 1.305908158532122e+17, 1.305908158655562e+17, 1.30590815877744e+17, 1.305908158899318e+17, 1.305908159021197e+17, 1.305908159143076e+17, 1.305908159266515e+17, 1.305908159388394e+17, 1.305908159510272e+17, 1.30590815963215e+17, 1.305908159754029e+17, 1.305908159877469e+17, 1.305908159999348e+17, 1.305908160121226e+17, 1.305908160243104e+17, 1.305908160364983e+17, 1.305908160488422e+17, 1.305908160610301e+17, 1.305908160732179e+17, 1.30590816085562e+17, 1.305908160977499e+17, 1.305908161099377e+17, 1.305908161221256e+17, 1.305908161344696e+17, 1.305908161466574e+17, 1.305908161588452e+17, 1.305908161710331e+17, 1.305908161832209e+17, 1.305908161954086e+17, 1.305908162077528e+17, 1.305908162199406e+17, 1.305908162321285e+17, 1.305908162443163e+17, 1.305908162565041e+17, 1.30590816268692e+17, 1.30590816281036e+17, 1.305908162932238e+17, 1.305908163054117e+17, 1.305908163175995e+17, 1.305908163297873e+17, 1.30590816341975e+17, 1.305908163543191e+17, 1.305908163665069e+17, 1.305908163786949e+17, 1.305908163908827e+17, 1.305908164030705e+17, 1.305908164152582e+17, 1.30590816427446e+17, 1.305908164397902e+17, 1.30590816451978e+17, 1.305908164641659e+17, 1.3059081647651e+17, 1.305908164885414e+17, 1.305908165008856e+17, 1.305908165130734e+17, 1.305908165252613e+17, 1.305908165374491e+17, 1.305908165496369e+17, 1.305908165619809e+17, 1.305908165741687e+17, 1.305908165863566e+17, 1.305908165985444e+17, 1.305908166107323e+17, 1.305908166230762e+17, 1.305908166352641e+17, 1.30590816647452e+17, 1.305908166596398e+17, 1.305908166718277e+17, 1.305908166840154e+17, 1.305908166963596e+17, 1.305908167085473e+17, 1.305908167207351e+17, 1.30590816732923e+17, 1.305908167452671e+17, 1.30590816757455e+17, 1.305908167696428e+17, 1.305908167818305e+17, 1.305908167940184e+17, 1.305908168062062e+17, 1.305908168185503e+17, 1.30590816830738e+17, 1.30590816842926e+17, 1.305908168551137e+17, 1.305908168673015e+17, 1.305908168794894e+17, 1.305908168918333e+17, 1.305908169040214e+17, 1.305908169162092e+17, 1.305908169283969e+17, 1.30590816940741e+17, 1.305908169527725e+17, 1.305908169651167e+17, 1.305908169773044e+17, 1.305908169894924e+17, 1.305908170016801e+17, 1.305908170140242e+17, 1.30590817026212e+17, 1.305908170383999e+17, 1.305908170507439e+17, 1.305908170629317e+17, 1.305908170751196e+17, 1.305908170873074e+17, 1.305908170994952e+17, 1.305908171118392e+17, 1.305908171240271e+17, 1.305908171362149e+17, 1.305908171484027e+17, 1.305908171605906e+17, 1.305908171727785e+17, 1.305908171851226e+17, 1.305908171973103e+17, 1.305908172094981e+17, 1.30590817221686e+17, 1.3059081723403e+17, 1.30590817246218e+17, 1.305908172584058e+17, 1.305908172705935e+17, 1.305908172827814e+17, 1.305908172951254e+17, 1.305908173073133e+17, 1.305908173195011e+17, 1.305908173318451e+17, 1.305908173440329e+17, 1.305908173562208e+17, 1.305908173684086e+17, 1.305908173805965e+17, 1.305908173927843e+17, 1.305908174051283e+17, 1.305908174173162e+17, 1.30590817429504e+17, 1.305908174416918e+17, 1.305908174538797e+17, 1.305908174662237e+17, 1.305908174784115e+17, 1.305908174905993e+17, 1.305908175027872e+17, 1.305908175149751e+17, 1.30590817527319e+17, 1.305908175395069e+17, 1.305908175516947e+17, 1.305908175638825e+17, 1.305908175762266e+17, 1.305908175884145e+17, 1.305908176006022e+17, 1.305908176129464e+17, 1.305908176251342e+17, 1.30590817637322e+17, 1.305908176496662e+17, 1.30590817661854e+17, 1.305908176740417e+17, 1.305908176862295e+17, 1.305908176984173e+17, 1.305908177106053e+17, 1.305908177227931e+17, 1.305908177351372e+17, 1.305908177473249e+17, 1.305908177595127e+17, 1.305908177718568e+17, 1.305908177840447e+17, 1.305908177962324e+17, 1.305908178084202e+17, 1.305908178206081e+17, 1.305908178329522e+17, 1.305908178451401e+17, 1.305908178573279e+17, 1.305908178695156e+17, 1.305908178817036e+17, 1.305908178938913e+17, 1.305908179062354e+17, 1.305908179184233e+17, 1.305908179306111e+17, 1.305908179427988e+17, 1.305908179549866e+17, 1.305908179673308e+17, 1.305908179795186e+17, 1.305908179917065e+17, 1.305908180038943e+17, 1.305908180160819e+17, 1.305908180282698e+17, 1.305908180404577e+17, 1.305908180528018e+17, 1.305908180649896e+17, 1.305908180771773e+17, 1.305908180893652e+17, 1.30590818101553e+17, 1.305908181138972e+17, 1.30590818126085e+17, 1.305908181382728e+17, 1.305908181504607e+17, 1.305908181628047e+17, 1.305908181749926e+17, 1.305908181871804e+17, 1.305908181993682e+17, 1.30590818211556e+17, 1.305908182239002e+17, 1.305908182360878e+17, 1.305908182482757e+17, 1.305908182604636e+17, 1.305908182728076e+17, 1.305908182849955e+17, 1.305908182971832e+17, 1.305908183093711e+17, 1.305908183215589e+17, 1.305908183337467e+17, 1.305908183460909e+17, 1.305908183582787e+17, 1.305908183704666e+17, 1.305908183826543e+17, 1.305908183948421e+17, 1.305908184071862e+17, 1.30590818419374e+17, 1.305908184315619e+17, 1.305908184437496e+17, 1.305908184559374e+17, 1.305908184681253e+17, 1.305908184804694e+17, 1.305908184926572e+17, 1.305908185048449e+17, 1.305908185170328e+17, 1.305908185292207e+17, 1.305908185415648e+17, 1.305908185537526e+17, 1.305908185659404e+17, 1.305908185781283e+17, 1.305908185904723e+17, 1.305908186026602e+17, 1.30590818614848e+17, 1.305908186270358e+17, 1.305908186392237e+17, 1.305908186515676e+17, 1.305908186637555e+17, 1.305908186759433e+17, 1.305908186881312e+17, 1.30590818700319e+17, 1.30590818712663e+17, 1.305908187248509e+17, 1.305908187370387e+17, 1.305908187492266e+17, 1.305908187614143e+17, 1.305908187737585e+17, 1.305908187859462e+17, 1.30590818798134e+17, 1.305908188104782e+17, 1.30590818822666e+17, 1.305908188348539e+17, 1.305908188470417e+17, 1.305908188592294e+17, 1.305908188715735e+17, 1.305908188837613e+17, 1.305908188959492e+17, 1.30590818908137e+17, 1.305908189203249e+17, 1.305908189325126e+17, 1.305908189448567e+17, 1.305908189570445e+17, 1.305908189692323e+17, 1.305908189814202e+17, 1.305908189936079e+17, 1.305908190057958e+17, 1.305908190181399e+17, 1.305908190303277e+17, 1.305908190425156e+17, 1.305908190547034e+17, 1.305908190668913e+17, 1.305908190792352e+17, 1.305908190914231e+17, 1.305908191036109e+17, 1.305908191157987e+17, 1.305908191281427e+17, 1.305908191403306e+17, 1.305908191525184e+17, 1.305908191648625e+17, 1.305908191770504e+17, 1.305908191892381e+17, 1.305908192014259e+17, 1.305908192136138e+17, 1.305908192258016e+17, 1.305908192381457e+17, 1.305908192503334e+17, 1.305908192625213e+17, 1.305908192747091e+17, 1.305908192868969e+17, 1.30590819299241e+17, 1.305908193114289e+17, 1.305908193236166e+17, 1.305908193358044e+17, 1.305908193479923e+17, 1.305908193601801e+17, 1.305908193725243e+17, 1.305908193847121e+17, 1.305908193968998e+17, 1.305908194090876e+17, 1.305908194212755e+17, 1.305908194336196e+17, 1.305908194458074e+17, 1.305908194579953e+17, 1.30590819470183e+17, 1.305908194823707e+17, 1.305908194945586e+17, 1.305908195069027e+17, 1.305908195190906e+17, 1.305908195312783e+17, 1.305908195436225e+17, 1.305908195558103e+17, 1.305908195679981e+17, 1.305908195801859e+17, 1.305908195925299e+17, 1.305908196047177e+17, 1.305908196169055e+17, 1.305908196290935e+17, 1.305908196414374e+17, 1.305908196536253e+17, 1.305908196658131e+17, 1.305908196781573e+17, 1.30590819690345e+17, 1.305908197025329e+17, 1.305908197147206e+17, 1.305908197269085e+17, 1.305908197392526e+17, 1.305908197514404e+17, 1.305908197636283e+17, 1.305908197758161e+17, 1.305908197880037e+17, 1.305908198003479e+17, 1.305908198125357e+17, 1.305908198247236e+17, 1.305908198369114e+17, 1.305908198492556e+17, 1.305908198614433e+17, 1.305908198736311e+17, 1.305908198858189e+17, 1.305908198980067e+17, 1.305908199103507e+17, 1.305908199225386e+17, 1.305908199347265e+17, 1.305908199469143e+17, 1.305908199591021e+17, 1.305908199714461e+17, 1.305908199836339e+17, 1.305908199958218e+17, 1.305908200080096e+17, 1.305908200201975e+17, 1.305908200323853e+17, 1.305908200447293e+17, 1.305908200569171e+17, 1.305908200691049e+17, 1.305908200812928e+17, 1.305908200934806e+17, 1.305908201056684e+17, 1.305908201180124e+17, 1.305908201302003e+17, 1.305908201423881e+17, 1.30590820154576e+17, 1.305908201669201e+17, 1.305908201791078e+17, 1.305908201912957e+17, 1.305908202034834e+17, 1.305908202156713e+17, 1.305908202278591e+17, 1.305908202402031e+17, 1.30590820252391e+17, 1.305908202645788e+17, 1.305908202769229e+17, 1.305908202891107e+17, 1.305908203012986e+17, 1.305908203134863e+17, 1.305908203256741e+17, 1.305908203380183e+17, 1.305908203502061e+17, 1.30590820362394e+17, 1.305908203745818e+17, 1.305908203869258e+17, 1.305908203991136e+17, 1.305908204113014e+17, 1.305908204234892e+17, 1.305908204356771e+17, 1.30590820447865e+17, 1.305908204602089e+17, 1.305908204723968e+17, 1.305908204845846e+17, 1.305908204967724e+17, 1.305908205089603e+17, 1.30590820521148e+17, 1.305908205334922e+17, 1.3059082054568e+17, 1.305908205578678e+17, 1.305908205700557e+17, 1.305908205823997e+17, 1.305908205945875e+17, 1.305908206067753e+17, 1.305908206189631e+17, 1.305908206313071e+17, 1.30590820643495e+17, 1.305908206556828e+17, 1.305908206678706e+17, 1.305908206800585e+17, 1.305908206922463e+17, 1.305908207045903e+17, 1.305908207167781e+17, 1.30590820728966e+17, 1.305908207411539e+17, 1.305908207533417e+17, 1.305908207656858e+17, 1.305908207778735e+17, 1.305908207900613e+17, 1.305908208022491e+17, 1.30590820814437e+17, 1.305908208266248e+17, 1.305908208388127e+17, 1.305908208511567e+17, 1.305908208633445e+17, 1.305908208755324e+17, 1.305908208877202e+17, 1.30590820899908e+17, 1.30590820912252e+17, 1.305908209244399e+17, 1.305908209366278e+17, 1.305908209488155e+17, 1.305908209610034e+17, 1.305908209733473e+17, 1.305908209855352e+17, 1.30590820997723e+17, 1.305908210100672e+17, 1.30590821022255e+17, 1.305908210344428e+17, 1.305908210466307e+17, 1.305908210588184e+17, 1.305908210711625e+17, 1.305908210833503e+17, 1.305908210955382e+17, 1.30590821107726e+17, 1.305908211199137e+17, 1.305908211322579e+17, 1.305908211444457e+17, 1.305908211566336e+17, 1.305908211688212e+17, 1.305908211811654e+17, 1.305908211933532e+17, 1.30590821205541e+17, 1.305908212177289e+17, 1.305908212299167e+17, 1.305908212422609e+17, 1.305908212544486e+17, 1.305908212666364e+17, 1.305908212789804e+17, 1.305908212911683e+17, 1.30590821303356e+17, 1.305908213155438e+17, 1.305908213277317e+17, 1.305908213399195e+17, 1.305908213522637e+17, 1.305908213644515e+17, 1.305908213766392e+17, 1.305908213888271e+17, 1.305908214010149e+17, 1.305908214132028e+17, 1.305908214255468e+17, 1.305908214377347e+17, 1.305908214499224e+17, 1.305908214622665e+17, 1.305908214744543e+17, 1.305908214866422e+17, 1.3059082149883e+17, 1.305908215110177e+17, 1.305908215233619e+17, 1.305908215355497e+17, 1.305908215477376e+17, 1.305908215599254e+17, 1.305908215722694e+17, 1.305908215803946e+17, 1.305908215925824e+17, 1.305908216047702e+17, 1.305908216169581e+17, 1.305908216291459e+17, 1.305908216413336e+17, 1.305908216536778e+17, 1.305908216658656e+17, 1.305908216780535e+17, 1.305908216902413e+17, 1.305908217024291e+17, 1.305908217146168e+17, 1.305908217269609e+17, 1.305908217391488e+17, 1.305908217513366e+17, 1.305908217635245e+17, 1.305908217757123e+17, 1.305908217880563e+17, 1.305908218002441e+17, 1.30590821812432e+17, 1.305908218246198e+17, 1.305908218368076e+17, 1.305908218491517e+17, 1.305908218613395e+17, 1.305908218735273e+17, 1.305908218857151e+17, 1.305908218979028e+17, 1.305908219100908e+17, 1.305908219222785e+17, 1.305908219344664e+17, 1.305908219466543e+17, 1.305908219589983e+17, 1.30590821971186e+17, 1.305908219833738e+17, 1.305908219914991e+17, 1.30590822003687e+17, 1.30590822016031e+17, 1.305908220282189e+17, 1.305908220404068e+17, 1.305908220525944e+17, 1.305908220647823e+17, 1.305908220771264e+17, 1.305908220893142e+17, 1.30590822101502e+17, 1.305908221136899e+17, 1.305908221258776e+17, 1.305908221382218e+17, 1.305908221504096e+17, 1.305908221625974e+17, 1.305908221749414e+17, 1.305908221869731e+17, 1.305908221993171e+17, 1.305908222115049e+17, 1.305908222236927e+17, 1.305908222360369e+17, 1.305908222482246e+17, 1.305908222604124e+17, 1.305908222726002e+17, 1.305908222849444e+17, 1.305908222971322e+17, 1.305908223093201e+17, 1.305908223215078e+17, 1.305908223336956e+17, 1.305908223460397e+17, 1.305908223582275e+17, 1.305908223705715e+17, 1.305908223827594e+17, 1.305908223949472e+17, 1.30590822407135e+17, 1.305908224194792e+17, 1.305908224316669e+17, 1.305908224438548e+17, 1.305908224561988e+17, 1.305908224683867e+17, 1.305908224805745e+17, 1.305908224927622e+17, 1.305908225049501e+17, 1.305908225172941e+17, 1.305908225294821e+17, 1.305908225416699e+17, 1.305908225538577e+17, 1.305908225660454e+17, 1.305908225782332e+17, 1.305908225904211e+17, 1.305908226026089e+17, 1.305908226149531e+17, 1.305908226271409e+17, 1.305908226393286e+17, 1.305908226515165e+17, 1.305908226596417e+17, 1.305908226719857e+17, 1.305908226841736e+17, 1.305908226963613e+17, 1.305908227085492e+17, 1.30590822720737e+17, 1.305908227288623e+17, 1.305908227410501e+17, 1.305908227533942e+17, 1.30590822765582e+17, 1.305908227777699e+17, 1.305908227899576e+17, 1.305908228021454e+17, 1.305908228143333e+17, 1.305908228266772e+17, 1.305908228388652e+17, 1.305908228510529e+17, 1.305908228632407e+17, 1.305908228755849e+17, 1.305908228877727e+17, 1.305908228999604e+17, 1.305908229121484e+17, 1.305908229243361e+17, 1.30590822936524e+17, 1.305908229488681e+17, 1.305908229610559e+17, 1.305908229732436e+17, 1.305908229855877e+17, 1.305908229977755e+17, 1.305908230099634e+17, 1.305908230221512e+17, 1.305908230343391e+17, 1.305908230466831e+17, 1.305908230588709e+17, 1.305908230710587e+17, 1.305908230832465e+17, 1.305908230954344e+17, 1.305908231077784e+17, 1.305908231199663e+17, 1.305908231321541e+17, 1.305908231441856e+17, 1.305908231563735e+17, 1.305908231687174e+17, 1.305908231809053e+17, 1.305908231930931e+17, 1.305908232052809e+17, 1.305908232174689e+17, 1.305908232298129e+17, 1.305908232420008e+17, 1.305908232541885e+17, 1.305908232663763e+17, 1.305908232785642e+17, 1.305908232909083e+17, 1.305908233030962e+17, 1.30590823315284e+17, 1.305908233274717e+17, 1.305908233398158e+17, 1.305908233520036e+17, 1.305908233641914e+17, 1.305908233763791e+17, 1.30590823388567e+17, 1.305908234007548e+17, 1.30590823413099e+17, 1.305908234252868e+17, 1.305908234374746e+17, 1.305908234496625e+17, 1.305908234618502e+17, 1.305908234741943e+17, 1.305908234863821e+17, 1.3059082349857e+17, 1.305908235107579e+17, 1.305908235229455e+17, 1.305908235351334e+17, 1.305908235473212e+17, 1.305908235596653e+17, 1.305908235718531e+17, 1.30590823584041e+17, 1.305908235962287e+17, 1.305908236084165e+17, 1.305908236206044e+17, 1.305908236327922e+17, 1.305908236451364e+17, 1.305908236573242e+17, 1.305908236695119e+17, 1.305908236816998e+17, 1.305908236938876e+17, 1.305908237062317e+17, 1.305908237184195e+17, 1.305908237306074e+17, 1.305908237427951e+17, 1.305908237549829e+17, 1.305908237671708e+17, 1.305908237795148e+17, 1.305908237917027e+17, 1.305908238038904e+17, 1.305908238160783e+17, 1.305908238282661e+17, 1.305908238406102e+17, 1.305908238527981e+17, 1.305908238649857e+17, 1.305908238771736e+17, 1.305908238893614e+17, 1.305908239015493e+17, 1.305908239138934e+17, 1.305908239260812e+17, 1.305908239382691e+17, 1.305908239506131e+17, 1.305908239628009e+17, 1.305908239749887e+17, 1.305908239871766e+17, 1.305908239993644e+17, 1.305908240115521e+17, 1.305908240238963e+17, 1.30590824036084e+17, 1.305908240482719e+17, 1.305908240604596e+17, 1.305908240726476e+17, 1.305908240849916e+17, 1.305908240971794e+17, 1.305908241093673e+17, 1.305908241215551e+17, 1.305908241337428e+17, 1.305908241460869e+17, 1.305908241582748e+17, 1.305908241704626e+17, 1.305908241826504e+17, 1.305908241948383e+17, 1.30590824207026e+17, 1.305908242193701e+17, 1.305908242315579e+17, 1.305908242437458e+17, 1.305908242560897e+17, 1.305908242682778e+17, 1.305908242804655e+17, 1.305908242926533e+17, 1.305908243049974e+17, 1.305908243171852e+17, 1.305908243293731e+17, 1.305908243415608e+17, 1.305908243537486e+17, 1.305908243660927e+17, 1.305908243782806e+17, 1.305908243904685e+17, 1.305908244026563e+17, 1.30590824414844e+17, 1.305908244270318e+17, 1.305908244393759e+17, 1.305908244515636e+17, 1.305908244637516e+17, 1.305908244759395e+17, 1.305908244882834e+17, 1.305908245004713e+17, 1.305908245126591e+17, 1.30590824524847e+17, 1.305908245371909e+17, 1.305908245493788e+17, 1.305908245615666e+17, 1.305908245737545e+17, 1.305908245860986e+17, 1.305908245982863e+17, 1.305908246104742e+17, 1.305908246226619e+17, 1.305908246348498e+17, 1.305908246470376e+17, 1.305908246592253e+17, 1.305908246715695e+17, 1.305908246837573e+17, 1.305908246959452e+17, 1.30590824708133e+17, 1.305908247203208e+17, 1.305908247326648e+17, 1.305908247448526e+17, 1.305908247570406e+17, 1.305908247692283e+17, 1.305908247814162e+17, 1.30590824793604e+17, 1.305908248057917e+17, 1.305908248181358e+17, 1.305908248303236e+17, 1.305908248426678e+17, 1.305908248548556e+17, 1.305908248670435e+17, 1.305908248792312e+17, 1.30590824891419e+17, 1.305908249037631e+17, 1.30590824915951e+17, 1.305908249281388e+17, 1.305908249403265e+17, 1.305908249526706e+17, 1.305908249648585e+17, 1.305908249770463e+17, 1.30590824989234e+17, 1.305908250015782e+17, 1.30590825013766e+17, 1.305908250259538e+17, 1.305908250382979e+17, 1.305908250504858e+17, 1.305908250626735e+17, 1.305908250748613e+17, 1.305908250870492e+17, 1.30590825099237e+17, 1.305908251115811e+17, 1.305908251237688e+17, 1.305908251359566e+17, 1.305908251481446e+17, 1.305908251603324e+17, 1.305908251725202e+17, 1.305908251848643e+17, 1.30590825197052e+17, 1.305908252092399e+17, 1.305908252214277e+17, 1.305908252336156e+17, 1.305908252458034e+17, 1.305908252581475e+17, 1.305908252703352e+17, 1.30590825282523e+17, 1.305908252947109e+17, 1.305908253068987e+17, 1.305908253190865e+17, 1.305908253312744e+17, 1.305908253436184e+17, 1.305908253558062e+17, 1.30590825367994e+17, 1.305908253801819e+17, 1.305908253923697e+17, 1.305908254045574e+17, 1.305908254169016e+17, 1.305908254290894e+17, 1.305908254412773e+17, 1.305908254536212e+17, 1.305908254658092e+17, 1.305908254779969e+17, 1.30590825490341e+17, 1.305908255025288e+17, 1.305908255147167e+17, 1.305908255269044e+17, 1.305908255390922e+17, 1.305908255512801e+17, 1.305908255636242e+17, 1.305908255758121e+17, 1.305908255879999e+17, 1.305908256001876e+17, 1.305908256123756e+17, 1.305908256245633e+17, 1.305908256367511e+17, 1.305908256490952e+17, 1.305908256611267e+17, 1.305908256733146e+17, 1.305908256856586e+17, 1.305908256978464e+17, 1.305908257101905e+17, 1.305908257223785e+17, 1.305908257345661e+17, 1.30590825746754e+17, 1.305908257589418e+17, 1.305908257711296e+17, 1.305908257834738e+17, 1.305908257956614e+17, 1.305908258078495e+17, 1.305908258200372e+17, 1.305908258323813e+17, 1.305908258445691e+17, 1.305908258567569e+17, 1.305908258689448e+17, 1.305908258811324e+17, 1.305908258933203e+17, 1.305908259056644e+17, 1.305908259178523e+17, 1.305908259300401e+17, 1.305908259423841e+17, 1.30590825954572e+17, 1.305908259667598e+17, 1.305908259789476e+17, 1.305908259911355e+17, 1.305908260034796e+17, 1.305908260156673e+17, 1.305908260278551e+17, 1.30590826040043e+17, 1.305908260522308e+17, 1.305908260644186e+17, 1.305908260766063e+17, 1.305908260889505e+17, 1.305908261011383e+17, 1.305908261133261e+17, 1.30590826125514e+17, 1.305908261377018e+17, 1.305908261498897e+17, 1.305908261620774e+17, 1.305908261744215e+17, 1.305908261866094e+17, 1.305908261987972e+17, 1.305908262109851e+17, 1.305908262231727e+17, 1.305908262353605e+17, 1.305908262475484e+17, 1.305908262598925e+17, 1.305908262720804e+17, 1.305908262842682e+17, 1.305908262964559e+17, 1.305908263086437e+17, 1.305908263209879e+17, 1.305908263331757e+17, 1.305908263453635e+17, 1.305908263575514e+17, 1.305908263698953e+17, 1.305908263820833e+17, 1.305908263942711e+17, 1.305908264064589e+17, 1.305908264186467e+17, 1.305908264309907e+17, 1.305908264431785e+17, 1.305908264553663e+17, 1.305908264677105e+17, 1.305908264798982e+17, 1.305908264920861e+17, 1.305908265042739e+17, 1.30590826516618e+17, 1.305908265288058e+17, 1.305908265409935e+17, 1.305908265531814e+17, 1.305908265653693e+17, 1.305908265775571e+17, 1.305908265899012e+17, 1.30590826602089e+17, 1.305908266142767e+17, 1.305908266264645e+17, 1.305908266386524e+17, 1.305908266508402e+17, 1.305908266631844e+17, 1.305908266753722e+17, 1.305908266875599e+17, 1.305908266997478e+17, 1.305908267119356e+17, 1.305908267241235e+17, 1.305908267364675e+17, 1.305908267486554e+17, 1.305908267608433e+17, 1.305908267730309e+17, 1.305908267852188e+17, 1.305908267974066e+17, 1.305908268097507e+17, 1.305908268219384e+17, 1.305908268341263e+17, 1.305908268463142e+17, 1.30590826858502e+17, 1.305908268708461e+17, 1.305908268830339e+17, 1.305908268952218e+17, 1.305908269074095e+17, 1.305908269195973e+17, 1.305908269317852e+17, 1.30590826943973e+17, 1.305908269563171e+17, 1.305908269685048e+17, 1.305908269806927e+17, 1.305908269928805e+17, 1.305908270050683e+17, 1.305908270172562e+17, 1.30590827029444e+17, 1.30590827041788e+17, 1.305908270539758e+17, 1.305908270661637e+17, 1.305908270783515e+17, 1.305908270905393e+17, 1.305908271027272e+17, 1.305908271150711e+17, 1.305908271272591e+17, 1.305908271394469e+17, 1.305908271516347e+17, 1.305908271638226e+17, 1.305908271761665e+17, 1.305908271883544e+17, 1.305908272005421e+17, 1.3059082721273e+17, 1.305908272249179e+17, 1.305908272371057e+17, 1.305908272494497e+17, 1.305908272616375e+17, 1.305908272738254e+17, 1.305908272860132e+17, 1.305908272983572e+17, 1.305908273105452e+17, 1.305908273227329e+17, 1.305908273349208e+17, 1.305908273471086e+17, 1.305908273594527e+17, 1.305908273716404e+17, 1.305908273838284e+17, 1.305908273961723e+17, 1.305908274083602e+17, 1.305908274207043e+17, 1.305908274328922e+17, 1.305908274450799e+17, 1.305908274572677e+17, 1.305908274694556e+17, 1.305908274817996e+17, 1.305908274939875e+17, 1.305908275061752e+17, 1.30590827518363e+17, 1.305908275305509e+17, 1.30590827542895e+17, 1.305908275550828e+17, 1.305908275672705e+17, 1.305908275794584e+17, 1.305908275918025e+17, 1.305908276039904e+17, 1.305908276161782e+17, 1.305908276285222e+17, 1.3059082764071e+17, 1.305908276528978e+17, 1.305908276650857e+17, 1.305908276774298e+17, 1.305908276896177e+17, 1.305908277019616e+17, 1.305908277141495e+17, 1.305908277263373e+17, 1.305908277385252e+17, 1.30590827750713e+17, 1.305908277588381e+17, 1.305908277669633e+17, 1.305908277750886e+17, 1.305908277833701e+17, 1.305908277914953e+17, 1.305908277996205e+17, 1.305908278077457e+17, 1.305908278158708e+17, 1.30590827823996e+17, 1.305908278321212e+17, 1.305908278402465e+17, 1.30590827848528e+17, 1.305908278566532e+17, 1.305908278647784e+17, 1.305908278769663e+17, 1.30590827889154e+17, 1.305908279013418e+17, 1.305908279135297e+17, 1.305908279258738e+17, 1.305908279380616e+17, 1.305908279502493e+17, 1.305908279624372e+17, 1.305908279746252e+17, 1.305908279869692e+17, 1.30590827999157e+17, 1.305908280113448e+17, 1.305908280235327e+17, 1.305908280357204e+17, 1.305908280479082e+17, 1.305908280602523e+17, 1.305908280724402e+17, 1.305908280847843e+17, 1.30590828096972e+17, 1.305908281091598e+17, 1.305908281213476e+17, 1.305908281335355e+17, 1.305908281457234e+17, 1.305908281580675e+17, 1.305908281702552e+17, 1.30590828182443e+17, 1.305908281946309e+17, 1.305908282068187e+17, 1.305908282190065e+17, 1.305908282313505e+17, 1.305908282435384e+17, 1.305908282557262e+17, 1.30590828267914e+17, 1.305908282801019e+17, 1.305908282924458e+17, 1.305908283046337e+17, 1.305908283168215e+17, 1.305908283290094e+17, 1.305908283411972e+17, 1.305908283535412e+17, 1.305908283657292e+17, 1.305908283779169e+17, 1.305908283901048e+17, 1.305908284022926e+17, 1.305908284144803e+17, 1.305908284266683e+17, 1.305908284390122e+17, 1.305908284512001e+17, 1.305908284633879e+17, 1.305908284755757e+17, 1.305908284877636e+17, 1.305908285001076e+17, 1.305908285122954e+17, 1.305908285244832e+17, 1.305908285366711e+17, 1.305908285488589e+17, 1.305908285612031e+17, 1.305908285733908e+17, 1.305908285857349e+17, 1.305908285979227e+17, 1.305908286101105e+17, 1.305908286222984e+17, 1.305908286344861e+17, 1.30590828646674e+17, 1.305908286588618e+17, 1.305908286712059e+17, 1.305908286832374e+17, 1.305908286954253e+17, 1.305908287077693e+17, 1.305908287199571e+17, 1.305908287323013e+17, 1.305908287444891e+17, 1.305908287566769e+17, 1.305908287688646e+17, 1.305908287810524e+17, 1.305908287932403e+17, 1.305908288054282e+17, 1.30590828817616e+17, 1.305908288299601e+17, 1.305908288421478e+17, 1.305908288543357e+17, 1.305908288665235e+17, 1.305908288787113e+17, 1.305908288908992e+17, 1.30590828903087e+17, 1.30590828915431e+17, 1.305908289274627e+17, 1.305908289398067e+17, 1.305908289519945e+17, 1.305908289641823e+17, 1.305908289765265e+17, 1.305908289887142e+17, 1.305908290009021e+17, 1.305908290130899e+17, 1.305908290252777e+17, 1.305908290374655e+17, 1.305908290498097e+17, 1.305908290619974e+17, 1.305908290741852e+17, 1.305908290863731e+17, 1.305908290985609e+17, 1.305908291107487e+17, 1.305908291230927e+17, 1.305908291352805e+17, 1.305908291474684e+17, 1.305908291596562e+17, 1.305908291720004e+17, 1.305908291841882e+17, 1.305908291963759e+17, 1.305908292085638e+17, 1.305908292207515e+17, 1.305908292329394e+17, 1.305908292452835e+17, 1.305908292574714e+17, 1.305908292698153e+17, 1.305908292820032e+17, 1.30590829294191e+17, 1.305908293063789e+17, 1.305908293185667e+17, 1.305908293309107e+17, 1.305908293430986e+17, 1.305908293552864e+17, 1.305908293674743e+17, 1.305908293796621e+17, 1.305908293918497e+17, 1.305908294041939e+17, 1.305908294163817e+17, 1.305908294285695e+17, 1.305908294407574e+17, 1.305908294529452e+17, 1.305908294652892e+17, 1.305908294774771e+17, 1.305908294896649e+17, 1.305908295018527e+17, 1.305908295140406e+17, 1.305908295262284e+17, 1.305908295384161e+17, 1.305908295507603e+17, 1.305908295629481e+17, 1.305908295751359e+17, 1.305908295873236e+17, 1.305908295995116e+17, 1.305908296116993e+17, 1.305908296240435e+17, 1.305908296362313e+17, 1.305908296484191e+17, 1.30590829660607e+17, 1.305908296727946e+17, 1.305908296851388e+17, 1.305908296973266e+17, 1.305908297095144e+17, 1.305908297218586e+17, 1.305908297340463e+17, 1.305908297462342e+17, 1.30590829758422e+17, 1.305908297706098e+17, 1.305908297827976e+17, 1.305908297951418e+17, 1.305908298073295e+17, 1.305908298195173e+17, 1.305908298317052e+17, 1.305908298438929e+17, 1.305908298560808e+17, 1.305908298684248e+17, 1.305908298806127e+17, 1.305908298928005e+17, 1.305908299049883e+17, 1.305908299171762e+17, 1.305908299295203e+17, 1.30590829941708e+17},
			             {1.305907699126172e+17, 1.305907699207424e+17, 1.305907699288677e+17, 1.305907699369929e+17, 1.305907699451181e+17, 1.305907699532433e+17, 1.305907699613684e+17, 1.305907699696499e+17, 1.305907699777751e+17, 1.305907699859003e+17, 1.305907699940256e+17, 1.305907700021508e+17, 1.30590770010276e+17, 1.305907700184013e+17, 1.305907700266828e+17, 1.305907700348079e+17, 1.305907700429332e+17, 1.305907700510583e+17, 1.305907700591836e+17, 1.305907700673088e+17, 1.30590770075434e+17, 1.305907700835592e+17, 1.305907700916844e+17, 1.305907700998095e+17, 1.305907701080911e+17, 1.305907701162163e+17, 1.305907701243415e+17, 1.305907701324667e+17, 1.305907701405919e+17, 1.305907701487172e+17, 1.305907701568424e+17, 1.305907701649676e+17, 1.305907701730929e+17, 1.30590770181218e+17, 1.305907701894995e+17, 1.305907701976248e+17, 1.3059077020575e+17, 1.305907702138752e+17, 1.305907702220004e+17, 1.305907702301256e+17, 1.305907702382508e+17, 1.305907702465322e+17, 1.305907702546575e+17, 1.305907702627827e+17, 1.305907702709079e+17, 1.305907702790331e+17, 1.305907702871583e+17, 1.305907702952835e+17, 1.305907703034088e+17, 1.30590770311534e+17, 1.305907703196591e+17, 1.305907703279406e+17, 1.305907703360658e+17, 1.305907703441911e+17, 1.305907703523164e+17, 1.305907703604416e+17, 1.305907703685668e+17, 1.30590770376692e+17, 1.305907703848172e+17, 1.305907703929423e+17, 1.305907704010675e+17, 1.30590770409349e+17, 1.305907704174742e+17, 1.305907704255995e+17, 1.305907704337247e+17, 1.3059077044185e+17, 1.30590770449975e+17, 1.305907704581004e+17, 1.305907704662255e+17, 1.30590770474507e+17, 1.305907704826322e+17, 1.305907704907575e+17, 1.305907704988827e+17, 1.305907705070079e+17, 1.305907705151332e+17, 1.305907705232584e+17, 1.305907705315398e+17, 1.30590770539665e+17, 1.305907705477902e+17, 1.305907705559154e+17, 1.305907705640406e+17, 1.305907705721658e+17, 1.305907705802909e+17, 1.305907705884163e+17, 1.305907705966977e+17, 1.305907706046668e+17, 1.305907706129482e+17, 1.305907706210734e+17, 1.305907706291986e+17, 1.305907706373238e+17, 1.305907706456052e+17, 1.305907706537306e+17, 1.305907706618557e+17, 1.305907706699809e+17, 1.305907706781062e+17, 1.305907706862314e+17, 1.305907706943566e+17, 1.305907707024818e+17, 1.305907707107633e+17, 1.305907707188886e+17, 1.305907707270136e+17, 1.305907707351388e+17, 1.305907707432641e+17, 1.305907707513893e+17, 1.305907707595145e+17, 1.305907707676398e+17, 1.30590770775765e+17, 1.305907707840465e+17, 1.305907707921716e+17, 1.305907708002968e+17, 1.305907708084221e+17, 1.305907708165473e+17, 1.305907708246725e+17, 1.305907708327978e+17, 1.30590770840923e+17, 1.305907708492045e+17, 1.305907708573297e+17, 1.305907708654548e+17, 1.3059077087358e+17, 1.305907708817052e+17, 1.305907708898304e+17, 1.305907708979557e+17, 1.305907709060809e+17, 1.305907709143624e+17, 1.305907709224876e+17, 1.305907709306127e+17, 1.30590770938738e+17, 1.305907709468632e+17, 1.305907709549884e+17, 1.305907709631137e+17, 1.305907709712389e+17, 1.305907709793641e+17, 1.305907709874893e+17, 1.305907709956145e+17, 1.305907710037398e+17, 1.305907710120212e+17, 1.305907710201464e+17, 1.305907710282716e+17, 1.305907710363968e+17, 1.30590771044522e+17, 1.305907710526473e+17, 1.305907710607725e+17, 1.305907710688977e+17, 1.305907710771791e+17, 1.305907710853044e+17, 1.305907710934296e+17, 1.305907711015548e+17, 1.3059077110968e+17, 1.305907711178053e+17, 1.305907711259305e+17, 1.30590771134212e+17, 1.305907711423372e+17, 1.305907711504623e+17, 1.305907711585876e+17, 1.305907711667128e+17, 1.305907711749943e+17, 1.305907711831195e+17, 1.305907711912447e+17, 1.305907711993699e+17, 1.30590771207495e+17, 1.305907712156202e+17, 1.305907712237455e+17, 1.305907712318707e+17, 1.305907712399959e+17, 1.305907712481212e+17, 1.305907712562464e+17, 1.305907712645279e+17, 1.305907712726531e+17, 1.305907712807784e+17, 1.305907712889036e+17, 1.305907712970287e+17, 1.305907713051539e+17, 1.305907713134354e+17, 1.305907713215607e+17, 1.305907713296859e+17, 1.305907713378111e+17, 1.305907713459363e+17, 1.305907713540614e+17, 1.305907713621866e+17, 1.305907713703118e+17, 1.305907713784371e+17, 1.305907713867185e+17, 1.305907713948438e+17, 1.305907714029691e+17, 1.305907714110943e+17, 1.305907714192195e+17, 1.305907714273446e+17, 1.3059077143547e+17, 1.305907714437513e+17, 1.305907714518766e+17, 1.305907714600018e+17, 1.30590771468127e+17, 1.305907714764084e+17, 1.305907714845338e+17, 1.305907714926589e+17, 1.305907715007841e+17, 1.305907715089093e+17, 1.305907715170345e+17, 1.305907715251597e+17, 1.30590771533285e+17, 1.305907715415665e+17, 1.305907715496916e+17, 1.305907715578168e+17, 1.30590771565942e+17, 1.305907715740673e+17, 1.305907715821925e+17, 1.305907715903177e+17, 1.305907715985992e+17, 1.305907716067244e+17, 1.305907716148497e+17, 1.305907716229748e+17, 1.305907716311e+17, 1.305907716392252e+17, 1.305907716473504e+17, 1.305907716554757e+17, 1.305907716637572e+17, 1.305907716718824e+17, 1.305907716800077e+17, 1.305907716881329e+17, 1.30590771696258e+17, 1.305907717045395e+17, 1.305907717126647e+17, 1.305907717207899e+17, 1.305907717289151e+17, 1.305907717370404e+17, 1.305907717453217e+17, 1.30590771753447e+17, 1.305907717615722e+17, 1.305907717696974e+17, 1.305907717778226e+17, 1.305907717859479e+17, 1.305907717940731e+17, 1.305907718021983e+17, 1.305907718104797e+17, 1.305907718186051e+17, 1.305907718267302e+17, 1.305907718348554e+17, 1.305907718431369e+17, 1.305907718512621e+17, 1.305907718593874e+17, 1.305907718675126e+17, 1.305907718756378e+17, 1.305907718837629e+17, 1.305907718918881e+17, 1.305907719000134e+17, 1.305907719082949e+17, 1.305907719164201e+17, 1.305907719245453e+17, 1.305907719326705e+17, 1.305907719407956e+17, 1.305907719489208e+17, 1.305907719570461e+17, 1.305907719651713e+17, 1.305907719734528e+17, 1.305907719815781e+17, 1.305907719897033e+17, 1.305907719978285e+17, 1.305907720059538e+17, 1.30590772014079e+17, 1.305907720222042e+17, 1.305907720303293e+17, 1.305907720386108e+17, 1.30590772046736e+17, 1.305907720548613e+17, 1.305907720629865e+17, 1.305907720711117e+17, 1.305907720792369e+17, 1.30590772087362e+17, 1.305907720954872e+17, 1.305907721037687e+17, 1.305907721118939e+17, 1.305907721200191e+17, 1.305907721281444e+17, 1.305907721362697e+17, 1.305907721443949e+17, 1.305907721525201e+17, 1.305907721606454e+17, 1.305907721687706e+17, 1.30590772177052e+17, 1.305907721851772e+17, 1.305907721933024e+17, 1.305907722014276e+17, 1.305907722097091e+17, 1.305907722178344e+17, 1.305907722259596e+17, 1.305907722340847e+17, 1.305907722422099e+17, 1.305907722503351e+17, 1.305907722584603e+17, 1.305907722667418e+17, 1.305907722748669e+17, 1.305907722829923e+17, 1.305907722911174e+17, 1.305907722992426e+17, 1.305907723073679e+17, 1.305907723154931e+17, 1.305907723236183e+17, 1.305907723317436e+17, 1.30590772340025e+17, 1.305907723481503e+17, 1.305907723562755e+17, 1.305907723644006e+17, 1.30590772372526e+17, 1.305907723806511e+17, 1.305907723887763e+17, 1.305907723969015e+17, 1.305907724050267e+17, 1.305907724133082e+17, 1.305907724214333e+17, 1.305907724295585e+17, 1.305907724376838e+17, 1.30590772445809e+17, 1.305907724539343e+17, 1.305907724620595e+17, 1.305907724701847e+17, 1.305907724784662e+17, 1.305907724865914e+17, 1.305907724947165e+17, 1.30590772502998e+17, 1.305907725111232e+17, 1.305907725192485e+17, 1.305907725273737e+17, 1.305907725354989e+17, 1.305907725436242e+17, 1.305907725517494e+17, 1.305907725600308e+17, 1.30590772568156e+17, 1.305907725762812e+17, 1.305907725844064e+17, 1.305907725925316e+17, 1.305907726006568e+17, 1.305907726087821e+17, 1.305907726169073e+17, 1.305907726251887e+17, 1.30590772633314e+17, 1.305907726414392e+17, 1.305907726495644e+17, 1.305907726576896e+17, 1.305907726658149e+17, 1.305907726739401e+17, 1.305907726820653e+17, 1.305907726903468e+17, 1.305907726984719e+17, 1.305907727065972e+17, 1.305907727147224e+17, 1.305907727228476e+17, 1.305907727309728e+17, 1.30590772739098e+17, 1.305907727472232e+17, 1.305907727553484e+17, 1.305907727634737e+17, 1.30590772771755e+17, 1.305907727798803e+17, 1.305907727880056e+17, 1.305907727961308e+17, 1.30590772804256e+17, 1.305907728125375e+17, 1.305907728205065e+17, 1.305907728287878e+17, 1.305907728369132e+17, 1.305907728450383e+17, 1.305907728531635e+17, 1.305907728612888e+17, 1.30590772869414e+17, 1.305907728775392e+17, 1.305907728856644e+17, 1.305907728937896e+17, 1.305907729019148e+17, 1.305907729101962e+17, 1.305907729183214e+17, 1.305907729264466e+17, 1.305907729345719e+17, 1.305907729428534e+17, 1.305907729509786e+17, 1.305907729591039e+17, 1.305907729672291e+17, 1.305907729753542e+17, 1.305907729834796e+17, 1.305907729916047e+17, 1.305907729997299e+17, 1.305907730078551e+17, 1.305907730159803e+17, 1.305907730241056e+17, 1.305907730323871e+17, 1.305907730405123e+17, 1.305907730486374e+17, 1.305907730567626e+17, 1.305907730648878e+17, 1.305907730730131e+17, 1.305907730811383e+17, 1.305907730894198e+17, 1.30590773097545e+17, 1.305907731056703e+17, 1.305907731137955e+17, 1.305907731219206e+17, 1.305907731300458e+17, 1.305907731381711e+17, 1.305907731464525e+17, 1.305907731545778e+17, 1.30590773162703e+17, 1.305907731708282e+17, 1.305907731789535e+17, 1.305907731870787e+17, 1.305907731952038e+17, 1.30590773203329e+17, 1.305907732114542e+17, 1.305907732195794e+17, 1.305907732278609e+17, 1.30590773235986e+17, 1.305907732441114e+17, 1.305907732522365e+17, 1.305907732603617e+17, 1.30590773268487e+17, 1.305907732766122e+17, 1.305907732847374e+17, 1.305907732930189e+17, 1.305907733011441e+17, 1.305907733092694e+17, 1.305907733173946e+17, 1.305907733255197e+17, 1.305907733336451e+17, 1.305907733417702e+17, 1.305907733500517e+17, 1.305907733580206e+17, 1.305907733663021e+17, 1.305907733744273e+17, 1.305907733825524e+17, 1.305907733906776e+17, 1.305907733988029e+17, 1.305907734070844e+17, 1.305907734150533e+17, 1.305907734231786e+17, 1.305907734314601e+17, 1.305907734395853e+17, 1.305907734477105e+17, 1.305907734558356e+17, 1.30590773463961e+17, 1.305907734722423e+17, 1.305907734803676e+17, 1.305907734884928e+17, 1.30590773496618e+17, 1.305907735047433e+17, 1.305907735128685e+17, 1.3059077352115e+17, 1.305907735292753e+17, 1.305907735374003e+17, 1.305907735455255e+17, 1.305907735536507e+17, 1.305907735617759e+17, 1.305907735700575e+17, 1.305907735781827e+17, 1.305907735863078e+17, 1.305907735944332e+17, 1.305907736027145e+17, 1.305907736108398e+17, 1.30590773618965e+17, 1.305907736270902e+17, 1.305907736352154e+17, 1.305907736433407e+17, 1.305907736514659e+17, 1.305907736595912e+17, 1.305907736678726e+17, 1.305907736759978e+17, 1.30590773684123e+17, 1.305907736922482e+17, 1.305907737003735e+17, 1.305907737084987e+17, 1.305907737166239e+17, 1.305907737247491e+17, 1.305907737328742e+17, 1.305907737411557e+17, 1.305907737492809e+17, 1.305907737574061e+17, 1.305907737655314e+17, 1.305907737736566e+17, 1.305907737817818e+17, 1.305907737900632e+17, 1.305907737981884e+17, 1.305907738063137e+17, 1.305907738144389e+17, 1.305907738225641e+17, 1.305907738306894e+17, 1.305907738388146e+17, 1.305907738469398e+17, 1.305907738550651e+17, 1.305907738633464e+17, 1.305907738714717e+17, 1.305907738795969e+17, 1.305907738877221e+17, 1.305907738960036e+17, 1.305907739041288e+17, 1.30590773912254e+17, 1.305907739203793e+17, 1.305907739285044e+17, 1.305907739366296e+17, 1.305907739447548e+17, 1.3059077395288e+17, 1.305907739611615e+17, 1.305907739692867e+17, 1.30590773977412e+17, 1.305907739855373e+17, 1.305907739936625e+17, 1.305907740017876e+17, 1.305907740099128e+17, 1.30590774018038e+17, 1.305907740263195e+17, 1.305907740344447e+17, 1.3059077404257e+17, 1.305907740506952e+17, 1.305907740588204e+17, 1.305907740669455e+17, 1.305907740750708e+17, 1.30590774083196e+17, 1.305907740914775e+17, 1.305907740996027e+17, 1.305907741077279e+17, 1.305907741158531e+17, 1.305907741241345e+17, 1.305907741322597e+17, 1.30590774140385e+17, 1.305907741485102e+17, 1.305907741566355e+17, 1.305907741647607e+17, 1.305907741728859e+17, 1.305907741811674e+17, 1.305907741892925e+17, 1.305907741974177e+17, 1.30590774205543e+17, 1.305907742136682e+17, 1.305907742217935e+17, 1.305907742300749e+17, 1.305907742382002e+17, 1.305907742463254e+17, 1.305907742544506e+17, 1.305907742625757e+17, 1.305907742707009e+17, 1.305907742788261e+17, 1.305907742869513e+17, 1.305907742950765e+17, 1.305907743032018e+17, 1.305907743113271e+17, 1.305907743196086e+17, 1.305907743277338e+17, 1.305907743358589e+17, 1.305907743439841e+17, 1.305907743521094e+17, 1.305907743602346e+17, 1.305907743683598e+17, 1.305907743766413e+17, 1.305907743847666e+17, 1.305907743928918e+17, 1.30590774401017e+17, 1.305907744091421e+17, 1.305907744172673e+17, 1.305907744253925e+17, 1.305907744335177e+17, 1.305907744417992e+17, 1.305907744499244e+17, 1.305907744580497e+17, 1.305907744661748e+17, 1.305907744743002e+17, 1.305907744825816e+17, 1.305907744907068e+17, 1.30590774498832e+17, 1.305907745069572e+17, 1.305907745150824e+17, 1.305907745232077e+17, 1.305907745313329e+17, 1.305907745394582e+17, 1.305907745475834e+17, 1.305907745557084e+17, 1.305907745638336e+17, 1.305907745719589e+17, 1.305907745800841e+17, 1.305907745883656e+17, 1.305907745964908e+17, 1.305907746046159e+17, 1.305907746127412e+17, 1.305907746208666e+17, 1.305907746289917e+17, 1.305907746371169e+17, 1.305907746453984e+17, 1.305907746535236e+17, 1.305907746616488e+17, 1.30590774669774e+17, 1.305907746778993e+17, 1.305907746861806e+17, 1.305907746943059e+17, 1.305907747024312e+17, 1.305907747105564e+17, 1.305907747186816e+17, 1.305907747268068e+17, 1.30590774734932e+17, 1.305907747430572e+17, 1.305907747511823e+17, 1.305907747593075e+17, 1.30590774767589e+17, 1.305907747757143e+17, 1.305907747838395e+17, 1.305907747919648e+17, 1.3059077480009e+17, 1.305907748082152e+17, 1.305907748163404e+17, 1.305907748244655e+17, 1.305907748325908e+17, 1.305907748408722e+17, 1.305907748489975e+17, 1.305907748571228e+17, 1.30590774865248e+17, 1.305907748733732e+17, 1.305907748814984e+17, 1.305907748896236e+17, 1.305907748977487e+17, 1.305907749060302e+17, 1.305907749141554e+17, 1.305907749222806e+17, 1.305907749304059e+17, 1.305907749385311e+17, 1.305907749466564e+17, 1.305907749549377e+17, 1.30590774963063e+17, 1.305907749711882e+17, 1.305907749793134e+17, 1.305907749875949e+17, 1.305907749957201e+17, 1.305907750038452e+17, 1.305907750119706e+17, 1.305907750200957e+17, 1.305907750282211e+17, 1.305907750363462e+17, 1.305907750446277e+17, 1.305907750527529e+17, 1.305907750608781e+17, 1.305907750690033e+17, 1.305907750771284e+17, 1.305907750852536e+17, 1.305907750933789e+17, 1.305907751015041e+17, 1.305907751096293e+17, 1.305907751177546e+17, 1.305907751258798e+17, 1.305907751341613e+17, 1.305907751422865e+17, 1.305907751504116e+17, 1.30590775158537e+17, 1.305907751666621e+17, 1.305907751747875e+17, 1.305907751829126e+17, 1.305907751911941e+17, 1.305907751993193e+17, 1.305907752074445e+17, 1.305907752155697e+17, 1.305907752236948e+17, 1.3059077523182e+17, 1.305907752399452e+17, 1.305907752480705e+17, 1.30590775256352e+17, 1.305907752644772e+17, 1.305907752726024e+17, 1.305907752807277e+17, 1.305907752888529e+17, 1.305907752971343e+17, 1.305907753052595e+17, 1.305907753133847e+17, 1.3059077532151e+17, 1.305907753296352e+17, 1.305907753377605e+17, 1.305907753458857e+17, 1.305907753541672e+17, 1.305907753622924e+17, 1.305907753704175e+17, 1.305907753785427e+17, 1.305907753866679e+17, 1.305907753947931e+17, 1.305907754029184e+17, 1.305907754111999e+17, 1.305907754193251e+17, 1.305907754274502e+17, 1.305907754355754e+17, 1.305907754437007e+17, 1.305907754518259e+17, 1.305907754599511e+17, 1.305907754680763e+17, 1.305907754762015e+17, 1.305907754844831e+17, 1.305907754926083e+17, 1.305907755007334e+17, 1.305907755088588e+17, 1.305907755169839e+17, 1.305907755251091e+17, 1.305907755332343e+17, 1.305907755413595e+17, 1.305907755494847e+17, 1.305907755577663e+17, 1.305907755658915e+17, 1.305907755740166e+17, 1.305907755821418e+17, 1.30590775590267e+17, 1.305907755983923e+17, 1.305907756065175e+17, 1.305907756146427e+17, 1.305907756229242e+17, 1.305907756310493e+17, 1.305907756391747e+17, 1.305907756472998e+17, 1.30590775655425e+17, 1.305907756635503e+17, 1.305907756716755e+17, 1.30590775679957e+17, 1.305907756880822e+17, 1.305907756962074e+17, 1.305907757043325e+17, 1.305907757124577e+17, 1.305907757207393e+17, 1.305907757288645e+17, 1.305907757369897e+17, 1.305907757451149e+17, 1.305907757532401e+17, 1.305907757613652e+17, 1.305907757694906e+17, 1.305907757776157e+17, 1.305907757858972e+17, 1.305907757940224e+17, 1.305907758021477e+17, 1.305907758102729e+17, 1.305907758183982e+17, 1.305907758265233e+17, 1.305907758346486e+17, 1.305907758427738e+17, 1.305907758508989e+17, 1.305907758591804e+17, 1.305907758673056e+17, 1.305907758754309e+17, 1.305907758835561e+17, 1.305907758916813e+17, 1.305907758998065e+17, 1.305907759079316e+17, 1.305907759160568e+17, 1.305907759241821e+17, 1.305907759323073e+17, 1.305907759404325e+17, 1.30590775948714e+17, 1.305907759568393e+17, 1.305907759649645e+17, 1.305907759730898e+17, 1.30590775981215e+17, 1.305907759893402e+17, 1.305907759974653e+17, 1.305907760055905e+17, 1.305907760137157e+17, 1.305907760218409e+17, 1.305907760301224e+17, 1.305907760382477e+17, 1.305907760463729e+17, 1.30590776054498e+17, 1.305907760626232e+17, 1.305907760707485e+17, 1.305907760788737e+17, 1.305907760869989e+17, 1.305907760951241e+17, 1.305907761034056e+17, 1.305907761115309e+17, 1.305907761196561e+17, 1.305907761277814e+17, 1.305907761359066e+17, 1.305907761440317e+17, 1.305907761521569e+17, 1.305907761602821e+17, 1.305907761684073e+17, 1.305907761765325e+17, 1.305907761846577e+17, 1.305907761929393e+17, 1.305907762010644e+17, 1.305907762091896e+17, 1.305907762173148e+17, 1.305907762254401e+17, 1.305907762335653e+17, 1.305907762416906e+17, 1.305907762498157e+17, 1.305907762580972e+17, 1.305907762662225e+17, 1.305907762743476e+17, 1.30590776282473e+17, 1.305907762905981e+17, 1.305907762987233e+17, 1.305907763068485e+17, 1.305907763149737e+17, 1.305907763230989e+17, 1.305907763312241e+17, 1.305907763395055e+17, 1.305907763476308e+17, 1.30590776355756e+17, 1.305907763638812e+17, 1.305907763720065e+17, 1.305907763801317e+17, 1.305907763882569e+17, 1.305907763963822e+17, 1.305907764046636e+17, 1.305907764127889e+17, 1.30590776420914e+17, 1.305907764290392e+17, 1.305907764371644e+17, 1.305907764452896e+17, 1.305907764534148e+17, 1.305907764616964e+17, 1.305907764698216e+17, 1.305907764779468e+17, 1.305907764860719e+17, 1.305907764941971e+17, 1.305907765023224e+17, 1.305907765104476e+17, 1.305907765185728e+17, 1.305907765266981e+17, 1.305907765349795e+17, 1.305907765431048e+17, 1.3059077655123e+17, 1.305907765593551e+17, 1.305907765674804e+17, 1.305907765756056e+17, 1.305907765837308e+17, 1.30590776591856e+17, 1.305907765999812e+17, 1.305907766081064e+17, 1.30590776616388e+17, 1.305907766245132e+17, 1.305907766326383e+17, 1.305907766407635e+17, 1.305907766488887e+17, 1.30590776657014e+17, 1.305907766651392e+17, 1.305907766734207e+17, 1.305907766815459e+17, 1.30590776689671e+17, 1.305907766979525e+17, 1.305907767060777e+17, 1.30590776714203e+17, 1.305907767223282e+17, 1.305907767304534e+17, 1.305907767385787e+17, 1.30590776746704e+17, 1.305907767549853e+17, 1.305907767631107e+17, 1.305907767712357e+17, 1.30590776779361e+17, 1.305907767874862e+17, 1.305907767956114e+17, 1.305907768037366e+17, 1.30590776812018e+17, 1.305907768201432e+17, 1.305907768282685e+17, 1.305907768363937e+17, 1.305907768446752e+17, 1.305907768528004e+17, 1.305907768609256e+17, 1.305907768690508e+17, 1.305907768771761e+17, 1.305907768853012e+17, 1.305907768934266e+17, 1.305907769015517e+17, 1.305907769096769e+17, 1.305907769179584e+17, 1.305907769260836e+17, 1.305907769342089e+17, 1.305907769423341e+17, 1.305907769504593e+17, 1.305907769585844e+17, 1.305907769668659e+17, 1.305907769749912e+17, 1.305907769831164e+17, 1.305907769912416e+17, 1.305907769993668e+17, 1.30590777007492e+17, 1.305907770156172e+17, 1.305907770238986e+17, 1.305907770320238e+17, 1.305907770401491e+17, 1.305907770482743e+17, 1.305907770563996e+17, 1.305907770645248e+17, 1.3059077707265e+17, 1.305907770807752e+17, 1.305907770889005e+17, 1.305907770970257e+17, 1.305907771051508e+17, 1.305907771134323e+17, 1.305907771215575e+17, 1.305907771296827e+17, 1.305907771378079e+17, 1.305907771459332e+17, 1.305907771540584e+17, 1.305907771621836e+17, 1.305907771703087e+17, 1.30590777178434e+17, 1.305907771867154e+17, 1.305907771948407e+17, 1.305907772029659e+17, 1.305907772110912e+17, 1.305907772192164e+17, 1.305907772274979e+17, 1.30590777235623e+17, 1.305907772437482e+17, 1.305907772518734e+17, 1.305907772599987e+17, 1.305907772681239e+17, 1.305907772764054e+17, 1.305907772845307e+17, 1.305907772926559e+17, 1.305907773007811e+17, 1.305907773089062e+17, 1.305907773170314e+17, 1.305907773251566e+17, 1.305907773334381e+17, 1.305907773415633e+17, 1.305907773496884e+17, 1.305907773578136e+17, 1.305907773659389e+17, 1.305907773740643e+17, 1.305907773821894e+17, 1.305907773903146e+17, 1.305907773984399e+17, 1.305907774065651e+17, 1.305907774146903e+17, 1.305907774229718e+17, 1.30590777431097e+17, 1.305907774392223e+17, 1.305907774473473e+17, 1.305907774554725e+17, 1.305907774635978e+17, 1.30590777471723e+17, 1.305907774798482e+17, 1.305907774879735e+17, 1.305907774962548e+17, 1.305907775043802e+17, 1.305907775125053e+17, 1.305907775206305e+17, 1.305907775287558e+17, 1.30590777536881e+17, 1.305907775450062e+17, 1.305907775531315e+17, 1.305907775612567e+17, 1.305907775695382e+17, 1.305907775776634e+17, 1.305907775857885e+17, 1.305907775939137e+17, 1.305907776020389e+17, 1.305907776101641e+17, 1.305907776182894e+17, 1.305907776264146e+17, 1.305907776345398e+17, 1.305907776428212e+17, 1.305907776509464e+17, 1.305907776590717e+17, 1.305907776671969e+17, 1.305907776753221e+17, 1.305907776834474e+17, 1.305907776917288e+17, 1.305907776998541e+17, 1.305907777079793e+17, 1.305907777161044e+17, 1.305907777242298e+17, 1.305907777323549e+17, 1.305907777404801e+17, 1.305907777486053e+17, 1.305907777567305e+17, 1.305907777648557e+17, 1.30590777772981e+17, 1.305907777811062e+17, 1.305907777892314e+17, 1.305907777975128e+17, 1.30590777805638e+17, 1.305907778137633e+17, 1.305907778218885e+17, 1.305907778300137e+17, 1.305907778382953e+17, 1.305907778462642e+17, 1.305907778543894e+17, 1.305907778626708e+17, 1.30590777870796e+17, 1.305907778789213e+17, 1.305907778870465e+17, 1.305907778951717e+17, 1.305907779032969e+17, 1.305907779114221e+17, 1.305907779195473e+17, 1.305907779276726e+17, 1.30590777935954e+17, 1.305907779440792e+17, 1.305907779522044e+17, 1.305907779604859e+17, 1.305907779686111e+17, 1.305907779767363e+17, 1.305907779848616e+17, 1.305907779929869e+17, 1.305907780011121e+17, 1.305907780092372e+17, 1.305907780173624e+17, 1.305907780254877e+17, 1.305907780336129e+17, 1.305907780418944e+17, 1.305907780500196e+17, 1.305907780581448e+17, 1.3059077806627e+17, 1.305907780743951e+17, 1.305907780825204e+17, 1.305907780906456e+17, 1.305907780987708e+17, 1.305907781068961e+17, 1.305907781150212e+17, 1.305907781231465e+17, 1.305907781312717e+17, 1.30590778139397e+17, 1.305907781475222e+17, 1.305907781558036e+17, 1.305907781639288e+17, 1.305907781720541e+17, 1.305907781801793e+17, 1.305907781884608e+17, 1.30590778196586e+17, 1.305907782047112e+17, 1.305907782128364e+17, 1.305907782209615e+17, 1.305907782290867e+17, 1.30590778237212e+17, 1.305907782453372e+17, 1.305907782534624e+17, 1.305907782615877e+17, 1.305907782697129e+17, 1.305907782779944e+17, 1.305907782861196e+17, 1.305907782942447e+17, 1.3059077830237e+17, 1.305907783104952e+17, 1.305907783186204e+17, 1.305907783267456e+17, 1.305907783350271e+17, 1.305907783431524e+17, 1.305907783512776e+17, 1.305907783594028e+17, 1.305907783675279e+17, 1.305907783756531e+17, 1.305907783837783e+17, 1.305907783919036e+17, 1.305907784000288e+17, 1.305907784083103e+17, 1.305907784164355e+17, 1.305907784245606e+17, 1.30590778432686e+17, 1.305907784408111e+17, 1.305907784489363e+17, 1.305907784570616e+17, 1.305907784651868e+17, 1.305907784734683e+17, 1.305907784815935e+17, 1.305907784897187e+17, 1.30590778497844e+17, 1.305907785059692e+17, 1.305907785140942e+17, 1.305907785222195e+17, 1.305907785303447e+17, 1.3059077853847e+17, 1.305907785465952e+17, 1.305907785547204e+17, 1.305907785630019e+17, 1.305907785709709e+17, 1.305907785792522e+17, 1.305907785873775e+17, 1.305907785955027e+17, 1.30590778603628e+17, 1.305907786117532e+17, 1.305907786198784e+17, 1.305907786280036e+17, 1.305907786362851e+17, 1.305907786444102e+17, 1.305907786525354e+17, 1.305907786606606e+17, 1.305907786687858e+17, 1.305907786769111e+17, 1.305907786850364e+17, 1.305907786931616e+17, 1.305907787012868e+17, 1.305907787095683e+17, 1.305907787176934e+17, 1.305907787258186e+17, 1.305907787339438e+17, 1.305907787420691e+17, 1.305907787501943e+17, 1.305907787584758e+17, 1.305907787666011e+17, 1.305907787747263e+17, 1.305907787828515e+17, 1.305907787909766e+17, 1.305907787992581e+17, 1.305907788073833e+17, 1.305907788155086e+17, 1.305907788236338e+17, 1.30590778831759e+17, 1.305907788398842e+17, 1.305907788480093e+17, 1.305907788561347e+17, 1.30590778864416e+17, 1.305907788725413e+17, 1.305907788806665e+17, 1.305907788887917e+17, 1.305907788969169e+17, 1.30590778905042e+17, 1.305907789131674e+17, 1.305907789212927e+17, 1.305907789294179e+17, 1.305907789376993e+17, 1.305907789458245e+17, 1.305907789539497e+17, 1.305907789620749e+17, 1.305907789702001e+17, 1.305907789784817e+17, 1.305907789866068e+17, 1.30590778994732e+17, 1.305907790028572e+17, 1.305907790109824e+17, 1.305907790192639e+17, 1.305907790272329e+17, 1.305907790355142e+17, 1.305907790434833e+17, 1.305907790517647e+17, 1.305907790598899e+17, 1.305907790680152e+17, 1.305907790761404e+17, 1.305907790842656e+17, 1.305907790923909e+17, 1.305907791005161e+17, 1.305907791086413e+17, 1.305907791167665e+17, 1.305907791248916e+17, 1.305907791330168e+17, 1.305907791412984e+17, 1.305907791494236e+17, 1.305907791575488e+17, 1.30590779165674e+17, 1.305907791737992e+17, 1.305907791819245e+17, 1.305907791900497e+17, 1.305907791981748e+17, 1.305907792063002e+17, 1.305907792145816e+17, 1.305907792227068e+17, 1.305907792308321e+17, 1.305907792389573e+17, 1.305907792470825e+17, 1.30590779255364e+17, 1.305907792634892e+17, 1.305907792716143e+17, 1.305907792797395e+17, 1.305907792878647e+17, 1.3059077929599e+17, 1.305907793041152e+17, 1.305907793122404e+17, 1.305907793203657e+17, 1.305907793284909e+17, 1.305907793367724e+17, 1.305907793448974e+17, 1.305907793530227e+17, 1.305907793611479e+17, 1.305907793692732e+17, 1.305907793773984e+17, 1.305907793856799e+17, 1.305907793938051e+17, 1.305907794019304e+17, 1.305907794100556e+17, 1.305907794181807e+17, 1.305907794263059e+17, 1.305907794344311e+17, 1.305907794427127e+17, 1.305907794508379e+17, 1.305907794589631e+17, 1.305907794670883e+17, 1.305907794752134e+17, 1.305907794833386e+17, 1.305907794914639e+17, 1.305907794995891e+17, 1.305907795078706e+17, 1.305907795159958e+17, 1.30590779524121e+17, 1.305907795322463e+17, 1.305907795403715e+17, 1.305907795484966e+17, 1.30590779556622e+17, 1.305907795647471e+17, 1.305907795728723e+17, 1.305907795809975e+17, 1.30590779589279e+17, 1.305907795974043e+17, 1.305907796055295e+17, 1.305907796136545e+17, 1.305907796217798e+17, 1.305907796300613e+17, 1.305907796381865e+17, 1.305907796463117e+17, 1.305907796544369e+17, 1.305907796625622e+17, 1.305907796706874e+17, 1.305907796788125e+17, 1.305907796870941e+17, 1.305907796952192e+17, 1.305907797033445e+17, 1.305907797114697e+17, 1.30590779719595e+17, 1.305907797277202e+17, 1.305907797360015e+17, 1.305907797441268e+17, 1.305907797522522e+17, 1.305907797603773e+17, 1.305907797685025e+17, 1.305907797766277e+17, 1.305907797847529e+17, 1.305907797928781e+17, 1.305907798010033e+17, 1.305907798092847e+17, 1.305907798174099e+17, 1.305907798255351e+17, 1.305907798336604e+17, 1.305907798417857e+17, 1.305907798499109e+17, 1.305907798580361e+17, 1.305907798663176e+17, 1.305907798742866e+17, 1.305907798825679e+17, 1.305907798906932e+17, 1.305907798988184e+17, 1.305907799069437e+17, 1.305907799152251e+17, 1.305907799233504e+17, 1.305907799314756e+17, 1.305907799396008e+17, 1.30590779947726e+17, 1.305907799558511e+17, 1.305907799639763e+17, 1.305907799722579e+17, 1.30590779980383e+17, 1.305907799885083e+17, 1.305907799966335e+17, 1.305907800047587e+17, 1.30590780012884e+17, 1.305907800210092e+17, 1.305907800291343e+17, 1.305907800372596e+17, 1.30590780045541e+17, 1.305907800536663e+17, 1.305907800617915e+17, 1.305907800699167e+17, 1.30590780078042e+17, 1.305907800861672e+17, 1.305907800942924e+17, 1.305907801025738e+17, 1.30590780110699e+17, 1.305907801188242e+17, 1.305907801269494e+17, 1.305907801350747e+17, 1.305907801431999e+17, 1.305907801513251e+17, 1.305907801594502e+17, 1.305907801675756e+17, 1.305907801758569e+17, 1.305907801839822e+17, 1.305907801921074e+17, 1.305907802002326e+17, 1.305907802083579e+17, 1.305907802164832e+17, 1.305907802246084e+17, 1.305907802327336e+17, 1.305907802408588e+17, 1.305907802489839e+17, 1.305907802571091e+17, 1.305907802653906e+17, 1.305907802735158e+17, 1.305907802816411e+17, 1.305907802897663e+17, 1.305907802978915e+17, 1.305907803060168e+17, 1.30590780314142e+17, 1.305907803224233e+17, 1.305907803305485e+17, 1.305907803386738e+17, 1.30590780346799e+17, 1.305907803550804e+17, 1.305907803632058e+17, 1.305907803713309e+17, 1.305907803794561e+17, 1.305907803875814e+17, 1.305907803955503e+17, 1.305907804038318e+17, 1.30590780411957e+17, 1.305907804200822e+17, 1.305907804283636e+17, 1.305907804364888e+17, 1.30590780444614e+17, 1.305907804527393e+17, 1.305907804608645e+17, 1.305907804689897e+17, 1.30590780477115e+17, 1.305907804852402e+17, 1.305907804935217e+17, 1.305907805016468e+17, 1.30590780509772e+17, 1.305907805178973e+17, 1.305907805260225e+17, 1.305907805341477e+17, 1.30590780542273e+17, 1.305907805503982e+17, 1.305907805586797e+17, 1.305907805668049e+17, 1.3059078057493e+17, 1.305907805830552e+17, 1.305907805911804e+17, 1.305907805993056e+17, 1.305907806074309e+17, 1.305907806155561e+17, 1.305907806236813e+17, 1.305907806318066e+17, 1.305907806400879e+17, 1.305907806482132e+17, 1.305907806563384e+17, 1.305907806644637e+17, 1.305907806725889e+17, 1.305907806807141e+17, 1.305907806888393e+17, 1.305907806969646e+17, 1.305907807050898e+17, 1.305907807133713e+17, 1.305907807214964e+17, 1.305907807296216e+17, 1.305907807377468e+17, 1.305907807458721e+17, 1.305907807541535e+17, 1.305907807622788e+17, 1.30590780770404e+17, 1.305907807785292e+17, 1.305907807866543e+17, 1.305907807947795e+17, 1.305907808029048e+17, 1.305907808111862e+17, 1.305907808193115e+17, 1.305907808272805e+17, 1.30590780835562e+17, 1.305907808436872e+17, 1.305907808518124e+17, 1.305907808599375e+17, 1.305907808680628e+17, 1.305907808763442e+17, 1.305907808844695e+17, 1.305907808925947e+17, 1.305907809007199e+17, 1.305907809088451e+17, 1.305907809169704e+17, 1.305907809250956e+17, 1.305907809332207e+17, 1.305907809413459e+17, 1.305907809496274e+17, 1.305907809577526e+17, 1.305907809658779e+17, 1.305907809740031e+17, 1.305907809821284e+17, 1.305907809902536e+17, 1.305907809983788e+17, 1.305907810065041e+17, 1.305907810146292e+17, 1.305907810229107e+17, 1.305907810310359e+17, 1.305907810391611e+17, 1.305907810472863e+17, 1.305907810554115e+17, 1.305907810635366e+17, 1.30590781071662e+17, 1.305907810797871e+17, 1.305907810880686e+17, 1.305907810961938e+17, 1.30590781104319e+17, 1.305907811124443e+17, 1.305907811205695e+17, 1.305907811286948e+17, 1.3059078113682e+17, 1.305907811449452e+17, 1.305907811532266e+17, 1.305907811613518e+17, 1.30590781169477e+17, 1.305907811776023e+17, 1.305907811857275e+17, 1.305907811938527e+17, 1.305907812019779e+17, 1.30590781210103e+17, 1.305907812183845e+17, 1.305907812265097e+17, 1.305907812346349e+17, 1.305907812427602e+17, 1.305907812508854e+17, 1.305907812591668e+17, 1.305907812671359e+17, 1.305907812752612e+17, 1.305907812833864e+17, 1.305907812916678e+17, 1.305907812996367e+17, 1.305907813079182e+17, 1.305907813160434e+17, 1.305907813241686e+17, 1.305907813322939e+17, 1.305907813405752e+17, 1.305907813485443e+17, 1.305907813568257e+17, 1.305907813649509e+17, 1.305907813730761e+17, 1.305907813812014e+17, 1.305907813893265e+17, 1.305907813974518e+17, 1.305907814057331e+17, 1.305907814138584e+17, 1.305907814219837e+17, 1.305907814301089e+17, 1.305907814382341e+17, 1.305907814463594e+17, 1.305907814546408e+17, 1.305907814627661e+17, 1.305907814708913e+17, 1.305907814790164e+17, 1.305907814871416e+17, 1.305907814952668e+17, 1.305907815033921e+17, 1.305907815116736e+17, 1.305907815197988e+17, 1.30590781527924e+17, 1.305907815360492e+17, 1.305907815441743e+17, 1.305907815522996e+17, 1.305907815604248e+17, 1.3059078156855e+17, 1.305907815766753e+17, 1.305907815849567e+17, 1.30590781593082e+17, 1.305907816012072e+17, 1.305907816093324e+17, 1.305907816174577e+17, 1.305907816255828e+17, 1.305907816338643e+17, 1.305907816419896e+17, 1.305907816501148e+17, 1.3059078165824e+17, 1.305907816663652e+17, 1.305907816744904e+17, 1.305907816826156e+17, 1.305907816907407e+17, 1.305907816988659e+17, 1.305907817071475e+17, 1.305907817152727e+17, 1.305907817233979e+17, 1.305907817315232e+17, 1.305907817396484e+17, 1.305907817477736e+17, 1.305907817558988e+17, 1.305907817641802e+17, 1.305907817723055e+17, 1.305907817804307e+17, 1.305907817885559e+17, 1.305907817966812e+17, 1.305907818048064e+17, 1.305907818129316e+17, 1.305907818210568e+17, 1.30590781829182e+17, 1.305907818373071e+17, 1.305907818455887e+17, 1.305907818537138e+17, 1.305907818618391e+17, 1.305907818699643e+17, 1.305907818780895e+17, 1.305907818862148e+17, 1.305907818943401e+17, 1.305907819024652e+17, 1.305907819107468e+17, 1.305907819188718e+17, 1.305907819269971e+17, 1.305907819351223e+17, 1.305907819432475e+17, 1.305907819513728e+17, 1.30590781959498e+17, 1.305907819676232e+17, 1.305907819759046e+17, 1.305907819840298e+17, 1.30590781992155e+17, 1.305907820002802e+17, 1.305907820084054e+17, 1.305907820165307e+17, 1.30590782024656e+17, 1.305907820329373e+17, 1.305907820410627e+17, 1.305907820491878e+17, 1.30590782057313e+17, 1.305907820654383e+17, 1.305907820737197e+17, 1.305907820816887e+17, 1.305907820899702e+17, 1.305907820980955e+17, 1.305907821062207e+17, 1.305907821143459e+17, 1.30590782122471e+17, 1.305907821305962e+17, 1.305907821388777e+17, 1.30590782147003e+17, 1.305907821551282e+17, 1.305907821632534e+17, 1.305907821713786e+17, 1.305907821795039e+17, 1.305907821876291e+17, 1.305907821959105e+17, 1.305907822040357e+17, 1.305907822121609e+17, 1.305907822202862e+17, 1.305907822284114e+17, 1.305907822365366e+17, 1.305907822446619e+17, 1.305907822527871e+17, 1.305907822609123e+17, 1.305907822691937e+17, 1.305907822773189e+17, 1.305907822854442e+17, 1.305907822935694e+17, 1.305907823016945e+17, 1.305907823099761e+17, 1.30590782317945e+17, 1.305907823262264e+17, 1.305907823343516e+17, 1.305907823424769e+17, 1.305907823507584e+17, 1.305907823588836e+17, 1.305907823670088e+17, 1.30590782375134e+17, 1.305907823832593e+17, 1.305907823913844e+17, 1.305907823995096e+17, 1.305907824076348e+17, 1.305907824159164e+17, 1.305907824240416e+17, 1.305907824321668e+17, 1.305907824402921e+17, 1.305907824484173e+17, 1.305907824565425e+17, 1.305907824646676e+17, 1.305907824729491e+17, 1.305907824810743e+17, 1.305907824891995e+17, 1.305907824974811e+17, 1.305907825056063e+17, 1.305907825137315e+17, 1.305907825218566e+17, 1.305907825299818e+17, 1.30590782538107e+17, 1.305907825462323e+17, 1.305907825543575e+17, 1.30590782562639e+17, 1.305907825707642e+17, 1.305907825788895e+17, 1.305907825870147e+17, 1.305907825951398e+17, 1.305907826032652e+17, 1.305907826113903e+17, 1.305907826195155e+17, 1.305907826276407e+17, 1.305907826359223e+17, 1.305907826440475e+17, 1.305907826521727e+17, 1.305907826602979e+17, 1.30590782668423e+17, 1.305907826765482e+17, 1.305907826846735e+17, 1.305907826927987e+17, 1.305907827010802e+17, 1.305907827092054e+17, 1.305907827173306e+17, 1.305907827254559e+17, 1.305907827335811e+17, 1.305907827417064e+17, 1.305907827498316e+17, 1.305907827579567e+17, 1.305907827660819e+17, 1.305907827742071e+17, 1.305907827824886e+17, 1.305907827906138e+17, 1.305907827987391e+17, 1.305907828068643e+17, 1.305907828149894e+17, 1.305907828231146e+17, 1.305907828312399e+17, 1.305907828393651e+17, 1.305907828474903e+17, 1.305907828557718e+17, 1.305907828638971e+17, 1.305907828720223e+17, 1.305907828801475e+17, 1.305907828882728e+17, 1.30590782896398e+17, 1.305907829045231e+17, 1.305907829126483e+17, 1.305907829207735e+17, 1.30590782929055e+17, 1.305907829371802e+17, 1.305907829453053e+17, 1.305907829534307e+17, 1.305907829615558e+17, 1.30590782969681e+17, 1.305907829778063e+17, 1.305907829859315e+17, 1.30590782994213e+17, 1.305907830023382e+17, 1.305907830104635e+17, 1.305907830187448e+17, 1.305907830268701e+17, 1.305907830349953e+17, 1.305907830431205e+17, 1.305907830512458e+17, 1.30590783059371e+17, 1.305907830674962e+17, 1.305907830756214e+17, 1.305907830837466e+17, 1.305907830920282e+17, 1.305907831001533e+17, 1.305907831082785e+17, 1.305907831164037e+17, 1.305907831245289e+17, 1.305907831326542e+17, 1.305907831407794e+17, 1.305907831489046e+17, 1.305907831570299e+17, 1.305907831651551e+17, 1.305907831734365e+17, 1.305907831815617e+17, 1.30590783189687e+17, 1.305907831978122e+17, 1.305907832059374e+17, 1.305907832140626e+17, 1.305907832221878e+17, 1.30590783230313e+17, 1.305907832384381e+17, 1.305907832467197e+17, 1.305907832546886e+17, 1.305907832629701e+17, 1.305907832710953e+17, 1.305907832792205e+17, 1.305907832873458e+17, 1.30590783295471e+17, 1.305907833035963e+17, 1.305907833117215e+17, 1.305907833200029e+17, 1.305907833281281e+17, 1.305907833362534e+17, 1.305907833443786e+17, 1.305907833525038e+17, 1.30590783360629e+17, 1.305907833687542e+17, 1.305907833768794e+17, 1.305907833851608e+17, 1.30590783393286e+17, 1.305907834014113e+17, 1.305907834095365e+17, 1.305907834176617e+17, 1.30590783425787e+17, 1.305907834339122e+17, 1.305907834421937e+17, 1.305907834503188e+17, 1.305907834584442e+17, 1.305907834665693e+17, 1.305907834746945e+17, 1.305907834828197e+17, 1.30590783490945e+17, 1.305907834990702e+17, 1.305907835071954e+17, 1.305907835154769e+17, 1.30590783523602e+17, 1.305907835317272e+17, 1.305907835398525e+17, 1.305907835479776e+17, 1.305907835561029e+17, 1.305907835642282e+17, 1.305907835723534e+17, 1.305907835806349e+17, 1.305907835887601e+17, 1.305907835968852e+17, 1.305907836050106e+17, 1.305907836131357e+17, 1.305907836212609e+17, 1.305907836293862e+17, 1.305907836375114e+17, 1.305907836456365e+17, 1.305907836537618e+17, 1.305907836620433e+17, 1.305907836701684e+17, 1.305907836782936e+17, 1.305907836864188e+17, 1.305907836945441e+17, 1.305907837026693e+17, 1.305907837107945e+17, 1.305907837189198e+17, 1.30590783727045e+17, 1.305907837351702e+17, 1.305907837432955e+17, 1.305907837514207e+17, 1.305907837597021e+17, 1.305907837678273e+17, 1.305907837759525e+17, 1.305907837840777e+17, 1.305907837922029e+17, 1.305907838003281e+17, 1.305907838084534e+17, 1.305907838165786e+17, 1.305907838247039e+17, 1.305907838328291e+17, 1.305907838411105e+17, 1.305907838492357e+17, 1.305907838573609e+17, 1.305907838654861e+17, 1.305907838736114e+17, 1.305907838817367e+17, 1.30590783890018e+17, 1.305907838979871e+17, 1.305907839062685e+17, 1.305907839143937e+17, 1.305907839225189e+17, 1.305907839306441e+17, 1.305907839387693e+17, 1.305907839468946e+17, 1.305907839550198e+17, 1.305907839633012e+17, 1.305907839714264e+17, 1.305907839795516e+17, 1.305907839876769e+17, 1.305907839958021e+17, 1.305907840039273e+17, 1.305907840120526e+17, 1.305907840203341e+17, 1.305907840284593e+17, 1.305907840365846e+17, 1.305907840447098e+17, 1.305907840528349e+17, 1.305907840609601e+17, 1.305907840692416e+17, 1.305907840773669e+17, 1.305907840854921e+17, 1.305907840936172e+17, 1.305907841017425e+17, 1.305907841098676e+17, 1.305907841179928e+17, 1.305907841261181e+17, 1.305907841342433e+17, 1.305907841425248e+17, 1.3059078415065e+17, 1.305907841587752e+17, 1.305907841669005e+17, 1.305907841750257e+17, 1.305907841831508e+17, 1.305907841912762e+17, 1.305907841994013e+17, 1.305907842075265e+17, 1.30590784215808e+17, 1.305907842239332e+17, 1.305907842320584e+17, 1.305907842401836e+17, 1.305907842484652e+17, 1.30590784256434e+17, 1.305907842645594e+17, 1.305907842726845e+17, 1.305907842808097e+17, 1.305907842889349e+17, 1.305907842972164e+17, 1.305907843053416e+17, 1.305907843134668e+17, 1.305907843215921e+17, 1.305907843297172e+17, 1.305907843378426e+17, 1.305907843459677e+17, 1.305907843540929e+17, 1.305907843622181e+17, 1.305907843704996e+17, 1.305907843786248e+17, 1.3059078438675e+17, 1.305907843948753e+17, 1.305907844030004e+17, 1.305907844111256e+17, 1.305907844192509e+17, 1.305907844273761e+17, 1.305907844355013e+17, 1.305907844437828e+17, 1.305907844519081e+17, 1.305907844600333e+17, 1.305907844681585e+17, 1.305907844762838e+17, 1.30590784484409e+17, 1.305907844925341e+17, 1.305907845006593e+17, 1.305907845087845e+17, 1.30590784517066e+17, 1.305907845251912e+17, 1.305907845333165e+17, 1.305907845414417e+17, 1.305907845495668e+17, 1.30590784557692e+17, 1.305907845658172e+17, 1.305907845739425e+17, 1.305907845820678e+17, 1.30590784590193e+17, 1.305907845984745e+17, 1.305907846065997e+17, 1.305907846147249e+17, 1.305907846228502e+17, 1.305907846309752e+17, 1.305907846392568e+17, 1.30590784647382e+17, 1.305907846555072e+17, 1.305907846636324e+17, 1.305907846717576e+17, 1.30590784680039e+17, 1.305907846881642e+17, 1.305907846962894e+17, 1.305907847044147e+17, 1.305907847125399e+17, 1.305907847206652e+17, 1.305907847287904e+17, 1.305907847369156e+17, 1.305907847450408e+17, 1.305907847533222e+17, 1.305907847614474e+17, 1.305907847695727e+17, 1.30590784777698e+17, 1.305907847858232e+17, 1.305907847939484e+17, 1.305907848020736e+17, 1.305907848101988e+17, 1.30590784818324e+17, 1.305907848264492e+17, 1.305907848347306e+17, 1.305907848428559e+17, 1.305907848509811e+17, 1.305907848591063e+17, 1.305907848672316e+17, 1.305907848753568e+17, 1.30590784883482e+17, 1.305907848916072e+17, 1.305907848997325e+17, 1.30590784908014e+17, 1.305907849161391e+17, 1.305907849242643e+17, 1.305907849323896e+17, 1.305907849405148e+17, 1.3059078494864e+17, 1.305907849567652e+17, 1.305907849650467e+17, 1.305907849731718e+17, 1.305907849812972e+17, 1.305907849894223e+17, 1.305907849975475e+17, 1.305907850056727e+17, 1.305907850137979e+17, 1.305907850219232e+17, 1.305907850300484e+17, 1.305907850381737e+17, 1.305907850464552e+17, 1.305907850545804e+17, 1.305907850627055e+17, 1.305907850708308e+17, 1.305907850789559e+17, 1.305907850870811e+17, 1.305907850952064e+17, 1.305907851033316e+17, 1.305907851114568e+17, 1.305907851197382e+17, 1.305907851278634e+17, 1.305907851359887e+17, 1.305907851442701e+17, 1.305907851523954e+17, 1.305907851605206e+17, 1.305907851686459e+17, 1.305907851767711e+17, 1.305907851847401e+17, 1.305907851930214e+17, 1.305907852011468e+17, 1.305907852092719e+17, 1.305907852173971e+17, 1.305907852255223e+17, 1.305907852338039e+17, 1.305907852419291e+17, 1.305907852500543e+17, 1.305907852581795e+17, 1.305907852663046e+17, 1.305907852744298e+17, 1.305907852827113e+17, 1.305907852908366e+17, 1.305907852989618e+17, 1.30590785307087e+17, 1.305907853152123e+17, 1.305907853233375e+17, 1.305907853314627e+17, 1.305907853397441e+17, 1.305907853478693e+17, 1.305907853559946e+17, 1.305907853641198e+17, 1.30590785372245e+17, 1.305907853803703e+17, 1.305907853884955e+17, 1.30590785396777e+17, 1.305907854047459e+17, 1.305907854130273e+17, 1.305907854211525e+17, 1.305907854292778e+17, 1.30590785437403e+17, 1.305907854455282e+17, 1.305907854536534e+17, 1.305907854619348e+17, 1.305907854700602e+17, 1.305907854781853e+17, 1.305907854863105e+17, 1.305907854944358e+17, 1.30590785502561e+17, 1.305907855108425e+17, 1.305907855189677e+17, 1.305907855270929e+17, 1.30590785535218e+17, 1.305907855433434e+17, 1.305907855514685e+17, 1.305907855595937e+17, 1.305907855677189e+17, 1.305907855760004e+17, 1.305907855841256e+17, 1.305907855922508e+17, 1.305907856003761e+17, 1.305907856085014e+17, 1.305907856166264e+17, 1.305907856247517e+17, 1.305907856330331e+17, 1.305907856411584e+17, 1.305907856492836e+17, 1.305907856574088e+17, 1.305907856655341e+17, 1.305907856736594e+17, 1.305907856819407e+17, 1.30590785690066e+17, 1.305907856981912e+17, 1.305907857063164e+17, 1.305907857145979e+17, 1.305907857227231e+17, 1.305907857308484e+17, 1.305907857389736e+17, 1.305907857470988e+17, 1.305907857552239e+17, 1.305907857633491e+17, 1.305907857716306e+17, 1.305907857797558e+17, 1.30590785787881e+17, 1.305907857960063e+17, 1.305907858041315e+17, 1.305907858122566e+17, 1.30590785820382e+17, 1.305907858285071e+17, 1.305907858367886e+17, 1.305907858449138e+17, 1.30590785853039e+17, 1.305907858611643e+17, 1.305907858692896e+17, 1.305907858775709e+17, 1.3059078588554e+17, 1.305907858938214e+17, 1.305907859019466e+17, 1.305907859100718e+17, 1.30590785918197e+17, 1.305907859263222e+17, 1.305907859346036e+17, 1.305907859427288e+17, 1.305907859508541e+17, 1.305907859589793e+17, 1.305907859671045e+17, 1.305907859752297e+17, 1.305907859835113e+17, 1.305907859916365e+17, 1.305907859997618e+17, 1.305907860078868e+17, 1.305907860160122e+17, 1.305907860241373e+17, 1.305907860322625e+17, 1.30590786040544e+17, 1.30590786048513e+17, 1.305907860567945e+17, 1.305907860649197e+17, 1.305907860730449e+17, 1.3059078608117e+17, 1.305907860894516e+17, 1.305907860975768e+17, 1.30590786105702e+17, 1.305907861138272e+17, 1.305907861219524e+17, 1.305907861300777e+17, 1.30590786138359e+17, 1.305907861464844e+17, 1.305907861546095e+17, 1.305907861627347e+17, 1.3059078617086e+17, 1.305907861789852e+17, 1.305907861871104e+17, 1.305907861952357e+17, 1.305907862033609e+17, 1.305907862114861e+17, 1.305907862196113e+17, 1.305907862277364e+17, 1.305907862358616e+17, 1.305907862441432e+17, 1.305907862522684e+17, 1.305907862603936e+17, 1.305907862685188e+17, 1.30590786276644e+17},
			             {1.30590786276644e+17, 1.305907862847693e+17, 1.305907862930506e+17, 1.305907863011759e+17, 1.305907863093012e+17, 1.305907863174264e+17, 1.305907863255516e+17, 1.305907863336769e+17, 1.30590786341802e+17, 1.305907863499273e+17, 1.305907863580525e+17, 1.30590786366334e+17, 1.305907863744591e+17, 1.305907863825843e+17, 1.305907863908659e+17, 1.305907863989911e+17, 1.305907864071163e+17, 1.305907864152415e+17, 1.305907864233667e+17, 1.305907864314918e+17, 1.305907864396172e+17, 1.305907864478986e+17, 1.305907864560238e+17, 1.30590786464149e+17, 1.305907864722743e+17, 1.305907864803995e+17, 1.305907864885247e+17, 1.3059078649665e+17, 1.305907865047752e+17, 1.305907865129004e+17, 1.305907865210255e+17, 1.305907865293071e+17, 1.305907865374323e+17, 1.305907865455575e+17, 1.305907865536827e+17, 1.305907865618079e+17, 1.305907865699331e+17, 1.305907865780584e+17, 1.305907865861836e+17, 1.305907865943087e+17, 1.305907866025902e+17, 1.305907866107154e+17, 1.305907866188407e+17, 1.305907866269659e+17, 1.305907866350911e+17, 1.305907866432164e+17, 1.305907866513416e+17, 1.30590786659623e+17, 1.305907866677482e+17, 1.305907866758734e+17, 1.305907866839987e+17, 1.305907866921239e+17, 1.305907867004054e+17, 1.305907867085306e+17, 1.305907867166557e+17, 1.305907867247809e+17, 1.305907867329061e+17, 1.305907867410313e+17, 1.305907867491566e+17, 1.305907867572819e+17, 1.305907867654071e+17, 1.305907867735323e+17, 1.305907867816575e+17, 1.305907867899389e+17, 1.305907867980641e+17, 1.305907868061894e+17, 1.305907868143146e+17, 1.305907868224398e+17, 1.30590786830565e+17, 1.305907868386902e+17, 1.305907868469718e+17, 1.30590786855097e+17, 1.305907868632221e+17, 1.305907868713473e+17, 1.305907868794725e+17, 1.305907868875978e+17, 1.30590786895723e+17, 1.305907869038482e+17, 1.305907869119735e+17, 1.305907869200987e+17, 1.305907869282239e+17, 1.305907869363492e+17, 1.305907869444744e+17, 1.305907869525996e+17, 1.30590786960881e+17, 1.305907869690062e+17, 1.305907869771314e+17, 1.305907869852566e+17, 1.305907869933818e+17, 1.305907870015071e+17, 1.305907870096324e+17, 1.305907870177576e+17, 1.305907870258828e+17, 1.305907870341642e+17, 1.305907870422894e+17, 1.305907870504146e+17, 1.305907870586961e+17, 1.305907870668214e+17, 1.305907870749466e+17, 1.305907870830717e+17, 1.305907870911971e+17, 1.305907870993222e+17, 1.305907871074474e+17, 1.305907871155726e+17, 1.305907871238541e+17, 1.305907871319794e+17, 1.305907871401046e+17, 1.305907871482296e+17, 1.305907871563549e+17, 1.305907871644801e+17, 1.305907871726053e+17, 1.305907871807306e+17, 1.305907871888558e+17, 1.305907871971373e+17, 1.305907872052626e+17, 1.305907872133878e+17, 1.30590787221513e+17, 1.305907872296381e+17, 1.305907872377633e+17, 1.305907872458886e+17, 1.305907872540138e+17, 1.30590787262139e+17, 1.305907872704205e+17, 1.305907872785457e+17, 1.305907872866708e+17, 1.305907872947962e+17, 1.305907873029213e+17, 1.305907873110465e+17, 1.305907873191718e+17, 1.30590787327297e+17, 1.305907873355785e+17, 1.305907873437037e+17, 1.305907873518289e+17, 1.305907873599542e+17, 1.305907873680794e+17, 1.305907873762045e+17, 1.305907873843299e+17, 1.30590787392455e+17, 1.305907874005802e+17, 1.305907874088617e+17, 1.305907874169869e+17, 1.305907874251121e+17, 1.305907874332372e+17, 1.305907874413624e+17, 1.305907874494877e+17, 1.305907874576131e+17, 1.305907874658944e+17, 1.305907874740197e+17, 1.305907874821449e+17, 1.305907874902701e+17, 1.305907874983953e+17, 1.305907875065206e+17, 1.305907875146458e+17, 1.305907875227711e+17, 1.305907875308963e+17, 1.305907875391777e+17, 1.305907875473029e+17, 1.305907875554281e+17, 1.305907875635533e+17, 1.305907875716785e+17, 1.305907875799601e+17, 1.305907875880852e+17, 1.305907875962103e+17, 1.305907876043356e+17, 1.305907876124608e+17, 1.30590787620586e+17, 1.305907876288675e+17, 1.305907876368365e+17, 1.30590787645118e+17, 1.305907876532433e+17, 1.305907876613684e+17, 1.305907876694936e+17, 1.305907876776188e+17, 1.30590787685744e+17, 1.305907876938693e+17, 1.305907877019945e+17, 1.30590787710276e+17, 1.305907877184012e+17, 1.305907877265263e+17, 1.305907877346515e+17, 1.305907877427767e+17, 1.30590787750902e+17, 1.305907877590272e+17, 1.305907877671525e+17, 1.305907877752777e+17, 1.305907877835592e+17, 1.305907877916844e+17, 1.305907877998095e+17, 1.305907878079348e+17, 1.3059078781606e+17, 1.305907878241852e+17, 1.305907878323105e+17, 1.305907878404357e+17, 1.305907878485609e+17, 1.305907878568424e+17, 1.305907878649676e+17, 1.305907878730927e+17, 1.305907878812179e+17, 1.305907878893432e+17, 1.305907878974684e+17, 1.305907879055937e+17, 1.305907879137189e+17, 1.305907879218441e+17, 1.305907879299693e+17, 1.305907879380945e+17, 1.305907879463759e+17, 1.305907879545012e+17, 1.305907879626264e+17, 1.305907879707517e+17, 1.305907879788769e+17, 1.305907879870021e+17, 1.305907879952836e+17, 1.305907880034088e+17, 1.30590788011534e+17, 1.305907880196591e+17, 1.305907880277843e+17, 1.305907880360659e+17, 1.305907880441911e+17, 1.305907880523163e+17, 1.305907880604415e+17, 1.305907880685667e+17, 1.30590788076692e+17, 1.305907880848173e+17, 1.305907880929425e+17, 1.305907881010676e+17, 1.305907881093491e+17, 1.305907881174743e+17, 1.305907881255995e+17, 1.305907881337247e+17, 1.3059078814185e+17, 1.305907881499752e+17, 1.305907881582566e+17, 1.30590788166382e+17, 1.30590788174507e+17, 1.305907881826322e+17, 1.305907881907574e+17, 1.305907881988827e+17, 1.305907882070079e+17, 1.305907882152893e+17, 1.305907882234145e+17, 1.305907882315398e+17, 1.30590788239665e+17, 1.305907882477902e+17, 1.305907882559155e+17, 1.305907882641969e+17, 1.30590788272166e+17, 1.305907882802912e+17, 1.305907882884164e+17, 1.305907882966979e+17, 1.30590788304823e+17, 1.305907883129482e+17, 1.305907883210734e+17, 1.305907883291986e+17, 1.305907883373238e+17, 1.305907883454491e+17, 1.305907883535744e+17, 1.305907883618557e+17, 1.305907883699811e+17, 1.305907883781062e+17, 1.305907883863876e+17, 1.305907883943566e+17, 1.305907884026381e+17, 1.305907884107634e+17, 1.305907884188886e+17, 1.305907884270138e+17, 1.305907884351391e+17, 1.305907884432643e+17, 1.305907884513894e+17, 1.305907884595146e+17, 1.305907884676398e+17, 1.305907884759214e+17, 1.305907884840466e+17, 1.305907884921718e+17, 1.30590788500297e+17, 1.305907885084221e+17, 1.305907885165473e+17, 1.305907885246726e+17, 1.305907885329541e+17, 1.305907885410793e+17, 1.305907885492045e+17, 1.305907885573298e+17, 1.30590788565455e+17, 1.305907885735802e+17, 1.305907885817053e+17, 1.305907885898307e+17, 1.305907885981121e+17, 1.305907886062373e+17, 1.305907886143626e+17, 1.305907886224877e+17, 1.305907886306129e+17, 1.30590788638738e+17, 1.305907886468634e+17, 1.305907886549885e+17, 1.305907886631139e+17, 1.305907886713952e+17, 1.305907886795205e+17, 1.305907886876457e+17, 1.305907886957709e+17, 1.305907887038962e+17, 1.305907887120214e+17, 1.305907887201466e+17, 1.30590788728428e+17, 1.305907887365532e+17, 1.305907887446785e+17, 1.305907887528037e+17, 1.305907887609289e+17, 1.305907887690541e+17, 1.305907887771793e+17, 1.305907887854609e+17, 1.30590788793586e+17, 1.305907888017112e+17, 1.305907888098364e+17, 1.305907888179616e+17, 1.305907888260869e+17, 1.305907888343683e+17, 1.305907888424936e+17, 1.305907888506188e+17, 1.305907888587441e+17, 1.305907888668692e+17, 1.305907888749944e+17, 1.305907888831197e+17, 1.305907888912449e+17, 1.305907888993701e+17, 1.305907889076516e+17, 1.305907889157769e+17, 1.305907889239021e+17, 1.305907889320273e+17, 1.305907889401524e+17, 1.305907889482776e+17, 1.305907889564028e+17, 1.305907889646843e+17, 1.305907889728095e+17, 1.305907889809348e+17, 1.3059078898906e+17, 1.305907889971852e+17, 1.305907890053103e+17, 1.305907890134356e+17, 1.305907890215608e+17, 1.305907890296861e+17, 1.305907890379676e+17, 1.305907890460928e+17, 1.30590789054218e+17, 1.305907890623433e+17, 1.305907890704684e+17, 1.305907890785935e+17, 1.305907890867187e+17, 1.305907890948439e+17, 1.305907891029692e+17, 1.305907891112507e+17, 1.305907891193759e+17, 1.305907891275012e+17, 1.305907891356264e+17, 1.305907891437516e+17, 1.305907891518769e+17, 1.30590789160002e+17, 1.305907891681272e+17, 1.305907891762525e+17, 1.305907891843777e+17, 1.305907891926592e+17, 1.305907892007844e+17, 1.305907892089096e+17, 1.30590789217191e+17, 1.305907892253164e+17, 1.305907892334415e+17, 1.305907892415667e+17, 1.305907892496919e+17, 1.305907892578171e+17, 1.305907892659423e+17, 1.305907892740675e+17, 1.305907892821928e+17, 1.305907892904742e+17, 1.305907892985994e+17, 1.305907893067247e+17, 1.305907893148499e+17, 1.305907893229751e+17, 1.305907893311003e+17, 1.305907893392256e+17, 1.305907893475071e+17, 1.305907893556323e+17, 1.305907893637576e+17, 1.305907893718828e+17, 1.305907893800079e+17, 1.305907893882894e+17, 1.305907893964146e+17, 1.305907894045398e+17, 1.30590789412665e+17, 1.305907894207903e+17, 1.305907894289155e+17, 1.305907894370406e+17, 1.305907894451658e+17, 1.30590789453291e+17, 1.305907894614163e+17, 1.305907894696977e+17, 1.305907894776667e+17, 1.305907894859483e+17, 1.305907894940735e+17, 1.305907895021987e+17, 1.305907895104801e+17, 1.305907895186053e+17, 1.305907895267306e+17, 1.305907895348558e+17, 1.30590789542981e+17, 1.305907895511062e+17, 1.305907895592314e+17, 1.305907895673565e+17, 1.305907895754819e+17, 1.305907895837632e+17, 1.305907895918885e+17, 1.305907896000137e+17, 1.30590789608139e+17, 1.305907896162642e+17, 1.305907896243894e+17, 1.305907896325146e+17, 1.305907896406399e+17, 1.305907896489212e+17, 1.305907896570465e+17, 1.305907896651717e+17, 1.30590789673297e+17, 1.305907896814222e+17, 1.305907896895474e+17, 1.305907896976726e+17, 1.30590789705954e+17, 1.305907897140792e+17, 1.305907897222044e+17, 1.305907897303297e+17, 1.305907897384549e+17, 1.305907897465801e+17, 1.305907897547054e+17, 1.305907897628306e+17, 1.305907897709558e+17, 1.30590789779081e+17, 1.305907897872063e+17, 1.305907897954877e+17, 1.305907898036129e+17, 1.305907898117381e+17, 1.305907898198634e+17, 1.305907898279886e+17, 1.305907898361138e+17, 1.30590789844239e+17, 1.305907898523642e+17, 1.305907898604893e+17, 1.305907898686147e+17, 1.305907898767398e+17, 1.305907898850213e+17, 1.305907898931465e+17, 1.305907899012717e+17, 1.30590789909397e+17, 1.305907899175222e+17, 1.305907899256475e+17, 1.305907899337727e+17, 1.305907899418979e+17, 1.305907899501793e+17, 1.305907899583046e+17, 1.305907899664297e+17, 1.305907899745549e+17, 1.305907899826802e+17, 1.305907899908054e+17, 1.305907899990868e+17, 1.30590790007212e+17, 1.305907900153372e+17, 1.305907900234625e+17, 1.305907900317439e+17, 1.305907900398692e+17, 1.305907900479944e+17, 1.305907900561197e+17, 1.305907900642449e+17, 1.3059079007237e+17, 1.305907900804952e+17, 1.305907900886205e+17, 1.305907900969019e+17, 1.305907901050272e+17, 1.305907901131525e+17, 1.305907901212777e+17, 1.305907901294029e+17, 1.305907901375281e+17, 1.305907901458095e+17, 1.305907901539347e+17, 1.305907901620599e+17, 1.305907901701851e+17, 1.305907901784667e+17, 1.305907901865919e+17, 1.305907901947171e+17, 1.305907902028422e+17, 1.305907902109674e+17, 1.305907902190927e+17, 1.305907902272179e+17, 1.305907902353431e+17, 1.305907902434684e+17, 1.305907902515936e+17, 1.305907902597188e+17, 1.305907902680003e+17, 1.305907902759693e+17, 1.305907902842508e+17, 1.305907902922196e+17, 1.305907903005011e+17, 1.305907903086263e+17, 1.305907903167516e+17, 1.305907903248768e+17, 1.305907903331583e+17, 1.305907903412835e+17, 1.305907903492524e+17, 1.305907903573777e+17, 1.30590790365503e+17, 1.305907903737843e+17, 1.305907903819096e+17, 1.305907903900348e+17, 1.3059079039816e+17, 1.305907904062853e+17, 1.305907904144104e+17, 1.305907904225356e+17, 1.305907904306609e+17, 1.30590790438786e+17, 1.305907904470675e+17, 1.305907904551927e+17, 1.305907904633179e+17, 1.305907904714432e+17, 1.305907904797245e+17, 1.305907904878499e+17, 1.305907904958189e+17, 1.305907905039441e+17, 1.305907905122255e+17, 1.305907905201946e+17, 1.305907905284759e+17, 1.305907905364449e+17, 1.305907905447264e+17, 1.305907905528516e+17, 1.305907905609768e+17, 1.30590790569102e+17, 1.305907905772271e+17, 1.305907905853524e+17, 1.305907905934776e+17, 1.305907906017591e+17, 1.305907906098844e+17, 1.305907906180096e+17, 1.305907906261348e+17, 1.305907906342601e+17, 1.305907906423853e+17, 1.305907906506668e+17, 1.305907906587919e+17, 1.305907906669171e+17, 1.305907906750423e+17, 1.305907906831676e+17, 1.305907906912928e+17, 1.30590790699418e+17, 1.305907907075432e+17, 1.305907907156684e+17, 1.3059079072395e+17, 1.305907907319188e+17, 1.30590790740044e+17, 1.305907907481693e+17, 1.305907907562945e+17, 1.30590790764576e+17, 1.305907907727012e+17, 1.305907907808264e+17, 1.305907907889517e+17, 1.305907907970769e+17, 1.305907908053583e+17, 1.305907908134836e+17, 1.305907908216088e+17, 1.30590790829734e+17, 1.305907908378592e+17, 1.305907908459844e+17, 1.305907908542659e+17, 1.30590790862391e+17, 1.305907908705162e+17, 1.305907908786415e+17, 1.305907908867667e+17, 1.305907908948919e+17, 1.305907909030172e+17, 1.305907909111424e+17, 1.305907909192676e+17, 1.305907909275491e+17, 1.305907909356742e+17, 1.305907909437996e+17, 1.305907909519247e+17, 1.305907909600499e+17, 1.305907909681752e+17, 1.305907909763004e+17, 1.305907909844256e+17, 1.305907909927071e+17, 1.305907910008323e+17, 1.305907910089574e+17, 1.305907910170826e+17, 1.305907910252078e+17, 1.305907910333331e+17, 1.305907910414583e+17, 1.305907910495835e+17, 1.30590791057865e+17, 1.305907910659903e+17, 1.305907910741155e+17, 1.305907910822408e+17, 1.305907910903658e+17, 1.305907910984911e+17, 1.305907911066163e+17, 1.305907911147415e+17, 1.305907911230231e+17, 1.305907911311483e+17, 1.305907911392735e+17, 1.305907911473987e+17, 1.305907911555238e+17, 1.30590791163649e+17, 1.305907911719306e+17, 1.305907911800558e+17, 1.30590791188181e+17, 1.305907911963062e+17, 1.305907912044314e+17, 1.305907912125567e+17, 1.30590791220838e+17, 1.305907912289633e+17, 1.305907912370885e+17, 1.305907912452137e+17, 1.30590791253339e+17, 1.305907912614643e+17, 1.305907912695895e+17, 1.305907912777147e+17, 1.305907912859962e+17, 1.305907912941213e+17, 1.305907913022465e+17, 1.305907913103717e+17, 1.305907913184969e+17, 1.305907913266222e+17, 1.305907913347474e+17, 1.305907913430289e+17, 1.30590791351154e+17, 1.305907913592792e+17, 1.305907913674045e+17, 1.305907913755297e+17, 1.305907913836549e+17, 1.305907913917802e+17, 1.305907913999054e+17, 1.305907914080306e+17, 1.305907914163121e+17, 1.305907914244372e+17, 1.305907914325626e+17, 1.305907914406877e+17, 1.305907914488129e+17, 1.305907914569381e+17, 1.305907914650633e+17, 1.305907914733449e+17, 1.305907914814701e+17, 1.305907914895953e+17, 1.305907914977204e+17, 1.305907915058458e+17, 1.305907915139709e+17, 1.305907915220961e+17, 1.305907915303776e+17, 1.305907915385028e+17, 1.30590791546628e+17, 1.305907915547532e+17, 1.305907915628785e+17, 1.305907915710038e+17, 1.30590791579129e+17, 1.305907915872541e+17, 1.305907915955356e+17, 1.305907916036608e+17, 1.305907916117861e+17, 1.305907916199113e+17, 1.305907916280365e+17, 1.305907916361617e+17, 1.305907916442868e+17, 1.30590791652412e+17, 1.305907916606935e+17, 1.305907916688187e+17, 1.30590791676944e+17, 1.305907916850692e+17, 1.305907916931945e+17, 1.305907917013197e+17, 1.30590791709445e+17, 1.305907917175702e+17, 1.305907917256954e+17, 1.305907917338205e+17, 1.30590791742102e+17, 1.305907917502273e+17, 1.305907917583524e+17, 1.305907917664776e+17, 1.305907917746029e+17, 1.305907917827281e+17, 1.305907917910095e+17, 1.305907917991347e+17, 1.305907918072599e+17, 1.305907918153852e+17, 1.305907918235104e+17, 1.305907918316356e+17, 1.305907918397609e+17, 1.305907918478861e+17, 1.305907918560113e+17, 1.305907918642927e+17, 1.305907918724179e+17, 1.305907918805432e+17, 1.305907918886684e+17, 1.305907918967936e+17, 1.305907919050752e+17, 1.305907919132003e+17, 1.305907919211692e+17, 1.305907919294508e+17, 1.305907919375759e+17, 1.305907919457011e+17, 1.305907919538264e+17, 1.305907919619516e+17, 1.305907919702331e+17, 1.305907919783583e+17, 1.305907919864835e+17, 1.305907919946086e+17, 1.30590792002734e+17, 1.305907920110154e+17, 1.305907920191406e+17, 1.305907920272658e+17, 1.305907920353911e+17, 1.305907920435163e+17, 1.305907920516415e+17, 1.305907920597668e+17, 1.305907920680481e+17, 1.305907920761734e+17, 1.305907920842986e+17, 1.305907920924238e+17, 1.30590792100549e+17, 1.305907921088305e+17, 1.305907921169558e+17, 1.305907921250808e+17, 1.305907921332061e+17, 1.305907921413313e+17, 1.305907921494566e+17, 1.305907921575818e+17, 1.30590792165707e+17, 1.305907921738322e+17, 1.305907921821137e+17, 1.30590792190239e+17, 1.305907921983642e+17, 1.305907922064893e+17, 1.305907922146147e+17, 1.305907922227398e+17, 1.30590792230865e+17, 1.305907922391465e+17, 1.305907922472717e+17, 1.305907922553969e+17, 1.305907922635222e+17, 1.305907922716472e+17, 1.305907922797725e+17, 1.305907922878977e+17, 1.305907922960229e+17, 1.305907923043044e+17, 1.305907923124296e+17, 1.305907923205549e+17, 1.305907923286802e+17, 1.305907923368054e+17, 1.305907923449306e+17, 1.305907923530557e+17, 1.305907923611809e+17, 1.305907923693062e+17, 1.305907923774314e+17, 1.305907923855566e+17, 1.305907923936818e+17, 1.305907924019633e+17, 1.305907924100884e+17, 1.305907924182138e+17, 1.305907924263389e+17, 1.305907924344641e+17, 1.305907924425894e+17, 1.305907924507146e+17, 1.305907924588398e+17, 1.305907924671213e+17, 1.305907924752465e+17, 1.305907924833718e+17, 1.30590792491497e+17, 1.305907924996221e+17, 1.305907925077475e+17, 1.305907925158726e+17, 1.305907925239978e+17, 1.30590792532123e+17, 1.305907925404045e+17, 1.305907925485297e+17, 1.305907925566548e+17, 1.3059079256478e+17, 1.305907925729053e+17, 1.305907925810307e+17, 1.305907925891557e+17, 1.30590792597281e+17, 1.305907926055624e+17, 1.305907926136877e+17, 1.305907926218129e+17, 1.305907926299382e+17, 1.305907926380634e+17, 1.305907926461887e+17, 1.305907926543137e+17, 1.305907926624389e+17, 1.305907926705641e+17, 1.305907926788457e+17, 1.305907926869709e+17, 1.305907926950961e+17, 1.305907927032212e+17, 1.305907927113466e+17, 1.305907927196279e+17, 1.305907927277532e+17, 1.305907927357222e+17, 1.305907927440036e+17, 1.305907927521289e+17, 1.305907927602541e+17, 1.305907927683794e+17, 1.305907927765046e+17, 1.30590792784786e+17, 1.305907927929112e+17, 1.305907928010364e+17, 1.305907928091616e+17, 1.305907928213495e+17, 1.305907928336936e+17, 1.305907928457252e+17, 1.305907928538504e+17, 1.305907928621318e+17, 1.30590792870257e+17, 1.305907928783823e+17, 1.305907928863512e+17, 1.305907928946327e+17, 1.305907929027579e+17, 1.305907929108831e+17, 1.305907929190083e+17, 1.305907929271336e+17, 1.305907929352586e+17, 1.305907929433839e+17, 1.305907929516654e+17, 1.305907929597906e+17, 1.305907929679159e+17, 1.305907929760411e+17, 1.305907929841663e+17, 1.305907929922916e+17, 1.305907930005729e+17, 1.305907930086982e+17, 1.305907930168236e+17, 1.305907930249487e+17, 1.305907930330739e+17, 1.30590793041199e+17, 1.305907930493242e+17, 1.305907930574495e+17, 1.305907930657309e+17, 1.305907930738561e+17, 1.305907930819814e+17, 1.305907930901066e+17, 1.305907930982318e+17, 1.305907931063571e+17, 1.305907931144823e+17, 1.305907931226075e+17, 1.305907931307327e+17, 1.305907931390141e+17, 1.305907931471395e+17, 1.305907931552646e+17, 1.305907931633898e+17, 1.30590793171515e+17, 1.305907931796402e+17, 1.305907931877654e+17, 1.305907931958907e+17, 1.305907932041722e+17, 1.305907932122973e+17, 1.305907932204225e+17, 1.305907932285477e+17, 1.305907932368292e+17, 1.305907932449544e+17, 1.305907932530797e+17, 1.30590793261205e+17, 1.305907932693302e+17},
			             {1.305907932693302e+17, 1.305907932774554e+17, 1.305907932857368e+17, 1.30590793293862e+17, 1.305907933019873e+17, 1.305907933101125e+17, 1.305907933182377e+17, 1.30590793326363e+17, 1.305907933344882e+17, 1.305907933426134e+17, 1.305907933507386e+17, 1.305907933588637e+17, 1.305907933671452e+17, 1.305907933752704e+17, 1.305907933833956e+17, 1.305907933915209e+17, 1.305907933996461e+17, 1.305907934077713e+17, 1.305907934158966e+17, 1.305907934240218e+17, 1.305907934323032e+17, 1.305907934404284e+17, 1.305907934485536e+17, 1.305907934566789e+17, 1.305907934649604e+17, 1.305907934730856e+17, 1.305907934812109e+17, 1.305907934893359e+17, 1.305907934974612e+17, 1.305907935055864e+17, 1.305907935138679e+17, 1.305907935219932e+17, 1.305907935301183e+17, 1.305907935382435e+17, 1.305907935463688e+17, 1.30590793554494e+17, 1.305907935626191e+17, 1.305907935707443e+17, 1.305907935788696e+17, 1.305907935869948e+17, 1.305907935952763e+17, 1.305907936034015e+17, 1.305907936115268e+17, 1.30590793619652e+17, 1.305907936277772e+17, 1.305907936359025e+17, 1.305907936440276e+17, 1.305907936521528e+17, 1.305907936604343e+17, 1.305907936685595e+17, 1.305907936766847e+17, 1.305907936848099e+17, 1.305907936930915e+17, 1.305907937010604e+17, 1.305907937093418e+17, 1.30590793717467e+17, 1.305907937255923e+17, 1.305907937337175e+17, 1.305907937418427e+17, 1.305907937501242e+17, 1.305907937582493e+17, 1.305907937663747e+17, 1.305907937744998e+17, 1.30590793782625e+17, 1.305907937907503e+17, 1.305907937988755e+17, 1.305907938070007e+17, 1.305907938152822e+17, 1.305907938234074e+17, 1.305907938315327e+17, 1.305907938396579e+17, 1.30590793847783e+17, 1.305907938559082e+17, 1.305907938640334e+17, 1.305907938721586e+17, 1.305907938804401e+17, 1.305907938885654e+17, 1.305907938966906e+17, 1.305907939048159e+17, 1.305907939129411e+17, 1.305907939210662e+17, 1.305907939291914e+17, 1.305907939373166e+17, 1.305907939454419e+17, 1.305907939537234e+17, 1.305907939618486e+17, 1.305907939699739e+17, 1.305907939780989e+17, 1.305907939862241e+17, 1.305907939943494e+17, 1.305907940024746e+17, 1.305907940105998e+17, 1.305907940187251e+17, 1.305907940268503e+17, 1.305907940351318e+17, 1.30590794043257e+17, 1.305907940513823e+17, 1.305907940595075e+17, 1.305907940676326e+17, 1.305907940757578e+17, 1.305907940838831e+17, 1.305907940920083e+17, 1.305907941001335e+17, 1.30590794108415e+17, 1.305907941165402e+17, 1.305907941246653e+17, 1.305907941327905e+17, 1.305907941409158e+17, 1.30590794149041e+17, 1.305907941571663e+17, 1.305907941652915e+17, 1.305907941734167e+17, 1.305907941816982e+17, 1.305907941898234e+17, 1.305907941979487e+17, 1.305907942060739e+17, 1.30590794214199e+17, 1.305907942223244e+17, 1.305907942304495e+17, 1.305907942385747e+17, 1.305907942466999e+17, 1.305907942548251e+17, 1.305907942629503e+17, 1.305907942712317e+17, 1.305907942793569e+17, 1.305907942874822e+17, 1.305907942956074e+17, 1.305907943037326e+17, 1.305907943118579e+17, 1.305907943199831e+17, 1.305907943281083e+17, 1.305907943362336e+17, 1.305907943443588e+17, 1.305907943526403e+17, 1.305907943607654e+17, 1.305907943688906e+17, 1.305907943770159e+17, 1.305907943851411e+17, 1.305907943932663e+17, 1.305907944013915e+17, 1.30590794409673e+17, 1.305907944177981e+17, 1.305907944259235e+17, 1.305907944340486e+17, 1.305907944423301e+17, 1.305907944504553e+17, 1.305907944585805e+17, 1.305907944667058e+17, 1.30590794474831e+17, 1.305907944829562e+17, 1.305907944912376e+17, 1.305907944993628e+17, 1.305907945074881e+17, 1.305907945156133e+17, 1.305907945237386e+17, 1.305907945318638e+17, 1.305907945401453e+17, 1.305907945482705e+17, 1.305907945563956e+17, 1.305907945645208e+17, 1.30590794572646e+17, 1.305907945807712e+17, 1.305907945888965e+17, 1.30590794597178e+17, 1.30590794605147e+17, 1.305907946134284e+17, 1.305907946215537e+17, 1.305907946296788e+17, 1.30590794637804e+17, 1.305907946460856e+17, 1.305907946542108e+17, 1.305907946621797e+17, 1.305907946704612e+17, 1.305907946785864e+17, 1.305907946867117e+17, 1.305907946948369e+17, 1.30590794702962e+17, 1.305907947110872e+17, 1.305907947192124e+17, 1.305907947273376e+17, 1.305907947354629e+17, 1.305907947435881e+17, 1.305907947517133e+17, 1.305907947598386e+17, 1.305907947679638e+17, 1.305907947762452e+17, 1.305907947843706e+17, 1.305907947924957e+17, 1.305907948006209e+17, 1.305907948087461e+17, 1.305907948168713e+17, 1.305907948249966e+17, 1.305907948331218e+17, 1.30590794841247e+17, 1.305907948493722e+17, 1.305907948576536e+17, 1.305907948657788e+17, 1.305907948739041e+17, 1.305907948820293e+17, 1.305907948901545e+17, 1.305907948982797e+17, 1.30590794906405e+17, 1.305907949145302e+17, 1.305907949228116e+17, 1.305907949309368e+17, 1.305907949390621e+17, 1.305907949473435e+17, 1.305907949554688e+17, 1.30590794963594e+17, 1.305907949717192e+17, 1.305907949798445e+17, 1.305907949879697e+17, 1.305907949960948e+17, 1.3059079500422e+17, 1.305907950123452e+17, 1.305907950204705e+17, 1.305907950285957e+17, 1.305907950368772e+17, 1.305907950450024e+17, 1.305907950531276e+17, 1.305907950612529e+17, 1.30590795069378e+17, 1.305907950775034e+17, 1.305907950857847e+17, 1.3059079509391e+17, 1.305907951020352e+17, 1.305907951101604e+17, 1.305907951182857e+17, 1.305907951264109e+17, 1.305907951345361e+17, 1.305907951428175e+17, 1.305907951509427e+17, 1.305907951590679e+17, 1.305907951671931e+17, 1.305907951753183e+17, 1.305907951834436e+17, 1.305907951915688e+17, 1.30590795199694e+17, 1.305907952078193e+17, 1.305907952159446e+17, 1.305907952242259e+17, 1.305907952323512e+17, 1.305907952404764e+17, 1.305907952486016e+17, 1.305907952567268e+17, 1.30590795264852e+17, 1.305907952729773e+17, 1.305907952811025e+17, 1.305907952893839e+17, 1.305907952975091e+17, 1.305907953056343e+17, 1.305907953137595e+17, 1.305907953218847e+17, 1.305907953301661e+17, 1.305907953381352e+17, 1.305907953464166e+17, 1.305907953545418e+17, 1.305907953626671e+17, 1.305907953707923e+17, 1.305907953789175e+17, 1.305907953870428e+17, 1.30590795395168e+17, 1.305907954034495e+17, 1.305907954115748e+17, 1.305907954196998e+17, 1.305907954278252e+17, 1.305907954359503e+17, 1.305907954440755e+17, 1.305907954522007e+17, 1.305907954604822e+17, 1.305907954686074e+17, 1.305907954767327e+17, 1.305907954848579e+17, 1.30590795492983e+17, 1.305907955011082e+17, 1.305907955092335e+17, 1.30590795517515e+17, 1.305907955256402e+17, 1.305907955337655e+17, 1.305907955418907e+17, 1.305907955500159e+17, 1.305907955581411e+17, 1.305907955662664e+17, 1.305907955743916e+17, 1.305907955825167e+17, 1.305907955906419e+17, 1.305907955989234e+17, 1.305907956070486e+17, 1.305907956151738e+17, 1.305907956232989e+17, 1.305907956314243e+17, 1.305907956395494e+17, 1.305907956476746e+17, 1.305907956557999e+17, 1.305907956639252e+17, 1.305907956720503e+17, 1.305907956801756e+17, 1.305907956883008e+17, 1.30590795696426e+17, 1.305907957047075e+17, 1.305907957128328e+17, 1.30590795720958e+17, 1.305907957290831e+17, 1.305907957372083e+17, 1.305907957453335e+17, 1.305907957534587e+17, 1.305907957617402e+17, 1.305907957698655e+17, 1.305907957779907e+17, 1.305907957861158e+17, 1.305907957942412e+17, 1.305907958023663e+17, 1.305907958104915e+17, 1.305907958186168e+17, 1.305907958268982e+17, 1.305907958350235e+17, 1.305907958431487e+17, 1.305907958512739e+17, 1.30590795859399e+17, 1.305907958675242e+17, 1.305907958756494e+17, 1.305907958837747e+17, 1.305907958918999e+17, 1.305907959000251e+17, 1.305907959083067e+17, 1.305907959164319e+17, 1.305907959245571e+17, 1.305907959326822e+17, 1.305907959408076e+17, 1.305907959489327e+17, 1.305907959570579e+17, 1.305907959651832e+17, 1.305907959734647e+17, 1.305907959815899e+17, 1.305907959897151e+17, 1.305907959978403e+17, 1.305907960059654e+17, 1.305907960140906e+17, 1.305907960222159e+17, 1.305907960303411e+17, 1.305907960386226e+17, 1.305907960467478e+17, 1.30590796054873e+17, 1.305907960629983e+17, 1.305907960712796e+17, 1.305907960794049e+17, 1.305907960875301e+17, 1.305907960956554e+17, 1.305907961037806e+17, 1.305907961119058e+17, 1.305907961200311e+17, 1.305907961283124e+17, 1.305907961364378e+17, 1.305907961445629e+17, 1.305907961526883e+17, 1.305907961608134e+17, 1.305907961689386e+17, 1.305907961770638e+17, 1.30590796185189e+17, 1.305907961934705e+17, 1.305907962015956e+17, 1.305907962097208e+17, 1.305907962178461e+17, 1.305907962259713e+17, 1.305907962340965e+17, 1.305907962422218e+17, 1.30590796250347e+17, 1.305907962584722e+17, 1.305907962667537e+17, 1.30590796274879e+17, 1.305907962830042e+17, 1.305907962911293e+17, 1.305907962992545e+17, 1.305907963073797e+17, 1.305907963155049e+17, 1.305907963237865e+17, 1.305907963319117e+17, 1.305907963400369e+17, 1.30590796348162e+17, 1.305907963564435e+17, 1.305907963645687e+17, 1.30590796372694e+17, 1.305907963808192e+17, 1.305907963889444e+17, 1.305907963970696e+17, 1.305907964051949e+17, 1.305907964133201e+17, 1.305907964214454e+17, 1.305907964297267e+17, 1.30590796437852e+17, 1.305907964459772e+17, 1.305907964541024e+17, 1.305907964622277e+17, 1.305907964701966e+17, 1.305907964784781e+17, 1.305907964866033e+17, 1.305907964947284e+17, 1.305907965030099e+17, 1.305907965111351e+17, 1.305907965192604e+17, 1.305907965273856e+17, 1.305907965355109e+17, 1.305907965436361e+17, 1.305907965517613e+17, 1.305907965598865e+17, 1.305907965680116e+17, 1.30590796576137e+17, 1.305907965842621e+17, 1.305907965923873e+17, 1.305907966005125e+17, 1.305907966087941e+17, 1.305907966169193e+17, 1.305907966250445e+17, 1.305907966331697e+17, 1.305907966412948e+17, 1.305907966494202e+17, 1.305907966577015e+17, 1.305907966658268e+17, 1.30590796673952e+17, 1.305907966820772e+17, 1.305907966902025e+17, 1.305907966983277e+17, 1.305907967064529e+17, 1.305907967147345e+17, 1.305907967228596e+17, 1.305907967309848e+17, 1.3059079673911e+17, 1.305907967472352e+17, 1.305907967553604e+17, 1.305907967634856e+17, 1.305907967716109e+17, 1.305907967798924e+17, 1.305907967880175e+17, 1.30590796796299e+17, 1.305907968044242e+17, 1.305907968125494e+17, 1.305907968206746e+17, 1.305907968287999e+17, 1.305907968369251e+17, 1.305907968450504e+17, 1.305907968533317e+17, 1.30590796861457e+17, 1.305907968695822e+17, 1.305907968777074e+17, 1.305907968858327e+17, 1.305907968939579e+17, 1.305907969020832e+17, 1.305907969102084e+17, 1.305907969184899e+17, 1.30590796926615e+17, 1.305907969347402e+17, 1.305907969428654e+17, 1.305907969509906e+17, 1.305907969591158e+17, 1.305907969672411e+17, 1.305907969753663e+17, 1.305907969834916e+17, 1.305907969916168e+17, 1.30590796999742e+17, 1.305907970078671e+17, 1.305907970159923e+17, 1.305907970242739e+17, 1.305907970323991e+17, 1.305907970405243e+17, 1.305907970486496e+17, 1.305907970567748e+17, 1.305907970649e+17, 1.305907970730252e+17, 1.305907970811503e+17, 1.305907970894318e+17, 1.30590797097557e+17, 1.305907971056822e+17, 1.305907971138075e+17, 1.305907971219327e+17, 1.305907971300579e+17, 1.305907971381832e+17, 1.305907971463084e+17, 1.305907971544335e+17, 1.305907971627151e+17, 1.305907971708403e+17},
			             {1.305907971708403e+17, 1.305907971789655e+17, 1.305907971870907e+17, 1.305907971952159e+17, 1.305907972033411e+17, 1.305907972114662e+17, 1.305907972197478e+17, 1.30590797227873e+17, 1.305907972359982e+17, 1.305907972441234e+17, 1.305907972522486e+17, 1.3059079726053e+17, 1.305907972684991e+17, 1.305907972766244e+17, 1.305907972847496e+17, 1.30590797293031e+17, 1.305907973011562e+17, 1.305907973092814e+17, 1.305907973174067e+17, 1.305907973255319e+17, 1.305907973378758e+17, 1.305907973500639e+17, 1.305907973622516e+17, 1.305907973745957e+17, 1.305907973866272e+17, 1.305907973989713e+17, 1.305907974111592e+17, 1.305907974192844e+17, 1.305907974274097e+17, 1.305907974358473e+17, 1.305907974477226e+17, 1.305907974599104e+17, 1.305907974722546e+17, 1.305907974844424e+17, 1.305907974966303e+17, 1.30590797508818e+17, 1.305907975169432e+17, 1.305907975252247e+17, 1.305907975374125e+17, 1.305907975455377e+17, 1.305907975578817e+17, 1.305907975700695e+17, 1.305907975822574e+17, 1.305907975903827e+17, 1.305907976025705e+17, 1.305907976106957e+17, 1.30590797618821e+17, 1.305907976271023e+17, 1.305907976352276e+17, 1.305907976474154e+17, 1.305907976555406e+17, 1.305907976677285e+17, 1.305907976758537e+17, 1.305907976839789e+17, 1.305907976963229e+17, 1.305907977044483e+17, 1.305907977125734e+17, 1.305907977247612e+17, 1.305907977328864e+17, 1.305907977410117e+17, 1.305907977491369e+17, 1.305907977572621e+17, 1.305907977655436e+17, 1.305907977777315e+17, 1.305907977899192e+17, 1.30590797802107e+17, 1.305907978103885e+17, 1.305907978185137e+17, 1.305907978307016e+17, 1.30590797838983e+17, 1.305907978511708e+17, 1.305907978633587e+17, 1.305907978755465e+17, 1.305907978836717e+17, 1.30590797891797e+17, 1.305907979041411e+17, 1.30590797916329e+17, 1.305907979244541e+17, 1.305907979366419e+17, 1.305907979447671e+17, 1.305907979569549e+17, 1.305907979652364e+17, 1.305907979733617e+17, 1.305907979814868e+17, 1.30590797989612e+17, 1.305907979977372e+17, 1.305907980100814e+17, 1.305907980222692e+17, 1.305907980303944e+17, 1.305907980385197e+17, 1.305907980507075e+17, 1.305907980588326e+17, 1.305907980710205e+17, 1.30590798079302e+17, 1.305907980914898e+17, 1.305907981036776e+17, 1.305907981158655e+17, 1.305907981280532e+17, 1.305907981403973e+17, 1.305907981525851e+17, 1.30590798164773e+17, 1.305907981769608e+17, 1.305907981893048e+17, 1.305907982014926e+17, 1.305907982136805e+17, 1.305907982258684e+17, 1.305907982380562e+17, 1.30590798250244e+17, 1.305907982624317e+17, 1.305907982747758e+17, 1.305907982869637e+17, 1.305907982991515e+17, 1.305907983113394e+17, 1.305907983235272e+17, 1.305907983358712e+17, 1.305907983480591e+17, 1.305907983602469e+17, 1.305907983724348e+17, 1.305907983846226e+17, 1.305907983968104e+17, 1.305907984089983e+17, 1.305907984213423e+17, 1.305907984335302e+17, 1.305907984457179e+17, 1.305907984579058e+17, 1.305907984700937e+17, 1.305907984824376e+17, 1.305907984946255e+17, 1.305907985068133e+17, 1.305907985191574e+17, 1.305907985313453e+17, 1.305907985435331e+17, 1.305907985557208e+17, 1.305907985679086e+17, 1.305907985802528e+17, 1.305907985924406e+17, 1.305907986046285e+17, 1.305907986168163e+17, 1.30590798629004e+17, 1.305907986411919e+17, 1.305907986533797e+17, 1.305907986655675e+17, 1.305907986777554e+17, 1.305907986899432e+17, 1.305907987021311e+17, 1.305907987143188e+17, 1.305907987266629e+17, 1.305907987388508e+17, 1.305907987510385e+17, 1.305907987633827e+17, 1.305907987755704e+17, 1.305907987877583e+17, 1.305907988001024e+17, 1.305907988122902e+17, 1.30590798824478e+17, 1.305907988366659e+17, 1.305907988488538e+17, 1.305907988611977e+17, 1.305907988733856e+17, 1.305907988857295e+17, 1.305907988979176e+17, 1.305907989101053e+17, 1.305907989224494e+17, 1.305907989346372e+17, 1.30590798946825e+17, 1.30590798959169e+17, 1.305907989713569e+17, 1.305907989835448e+17, 1.305907989957325e+17, 1.305907990079204e+17, 1.305907990201083e+17, 1.305907990322961e+17, 1.30590799044484e+17, 1.305907990566717e+17, 1.305907990688595e+17, 1.305907990812036e+17, 1.305907990933914e+17, 1.305907991055793e+17, 1.30590799117767e+17, 1.305907991299549e+17, 1.30590799142299e+17, 1.305907991544868e+17, 1.30590799162612e+17, 1.305907991747999e+17, 1.305907991830813e+17, 1.305907991952691e+17, 1.30590799207457e+17, 1.305907992196448e+17, 1.305907992318326e+17, 1.305907992440205e+17, 1.305907992562083e+17, 1.305907992685523e+17, 1.305907992807402e+17, 1.30590799292928e+17, 1.305907993051159e+17, 1.3059079931746e+17, 1.305907993296477e+17, 1.305907993418355e+17, 1.305907993540234e+17, 1.305907993662112e+17, 1.305907993785553e+17, 1.305907993866806e+17, 1.305907993988684e+17, 1.305907994110561e+17, 1.30590799423244e+17, 1.305907994354318e+17, 1.305907994476196e+17, 1.305907994598075e+17, 1.305907994721516e+17, 1.305907994843395e+17, 1.305907994965272e+17, 1.30590799508715e+17, 1.305907995209029e+17, 1.305907995330907e+17, 1.305907995454348e+17, 1.305907995576225e+17, 1.305907995698104e+17, 1.305907995821544e+17, 1.305907995943423e+17, 1.3059079960653e+17, 1.305907996187178e+17, 1.30590799631062e+17, 1.305907996432498e+17, 1.305907996554377e+17, 1.305907996676255e+17, 1.305907996799697e+17, 1.305907996921573e+17, 1.305907997043452e+17, 1.305907997165331e+17, 1.305907997288771e+17, 1.30590799741065e+17, 1.30590799753409e+17, 1.305907997655968e+17, 1.305907997777847e+17, 1.305907997901288e+17, 1.305907998023165e+17, 1.305907998145044e+17, 1.305907998266922e+17, 1.305907998390363e+17, 1.305907998512242e+17, 1.30590799863412e+17, 1.305907998755999e+17, 1.305907998879438e+17, 1.305907999001317e+17, 1.305907999123195e+17, 1.305907999245073e+17, 1.305907999366952e+17, 1.305907999488829e+17, 1.30590799961227e+17, 1.305907999734149e+17, 1.305907999856027e+17, 1.305907999977905e+17, 1.305908000099782e+17, 1.305908000223224e+17, 1.305908000345102e+17, 1.305908000466981e+17, 1.305908000588859e+17, 1.305908000710737e+17, 1.305908000834179e+17, 1.305908000956056e+17, 1.305908001077935e+17, 1.305908001199813e+17, 1.305908001323254e+17, 1.305908001445133e+17, 1.305908001567011e+17, 1.305908001688888e+17, 1.305908001812329e+17, 1.305908001934207e+17, 1.305908002056086e+17, 1.305908002177964e+17, 1.305908002301404e+17, 1.305908002423283e+17, 1.305908002545161e+17, 1.305908002667039e+17, 1.305908002788918e+17, 1.305908002912358e+17, 1.305908003034237e+17, 1.305908003156115e+17, 1.305908003279556e+17, 1.305908003401435e+17, 1.305908003523313e+17, 1.30590800364519e+17, 1.30590800376863e+17, 1.30590800389051e+17, 1.305908004012388e+17, 1.305908004134266e+17, 1.305908004256145e+17, 1.305908004378022e+17, 1.3059080044999e+17, 1.305908004623341e+17, 1.30590800474522e+17, 1.305908004867098e+17, 1.305908004988975e+17, 1.305908005110854e+17, 1.305908005234295e+17, 1.305908005356174e+17, 1.305908005478052e+17, 1.30590800559993e+17, 1.305908005721809e+17, 1.305908005843686e+17, 1.305908005967128e+17, 1.305908006089006e+17, 1.305908006210884e+17, 1.305908006332762e+17, 1.305908006454641e+17, 1.305908006576518e+17, 1.305908006698397e+17, 1.305908006821838e+17, 1.305908006943715e+17, 1.305908007065594e+17, 1.305908007187473e+17, 1.30590800730935e+17, 1.305908007431228e+17, 1.305908007554669e+17, 1.305908007676548e+17, 1.305908007798427e+17, 1.305908007920303e+17, 1.305908008042182e+17, 1.305908008165623e+17, 1.305908008287501e+17, 1.30590800840938e+17, 1.305908008531258e+17, 1.3059080086547e+17, 1.305908008776577e+17, 1.305908008898455e+17, 1.305908009020334e+17, 1.305908009143775e+17, 1.305908009265652e+17, 1.30590800938753e+17, 1.305908009509409e+17, 1.305908009631287e+17, 1.305908009754728e+17, 1.305908009876605e+17, 1.305908009998484e+17, 1.305908010120364e+17, 1.305908010242241e+17, 1.305908010364119e+17, 1.305908010485997e+17, 1.305908010609439e+17, 1.305908010731316e+17, 1.305908010853194e+17, 1.305908010975073e+17, 1.305908011096951e+17, 1.305908011220393e+17, 1.305908011342271e+17, 1.305908011464148e+17, 1.305908011586028e+17, 1.305908011707905e+17, 1.305908011829783e+17, 1.305908011951662e+17, 1.305908012075103e+17, 1.30590801219698e+17, 1.305908012320421e+17, 1.3059080124423e+17, 1.305908012564177e+17, 1.305908012686056e+17, 1.305908012807935e+17, 1.305908012931375e+17, 1.305908013053253e+17, 1.305908013175131e+17, 1.30590801329701e+17, 1.305908013418888e+17, 1.305908013540765e+17, 1.305908013664207e+17, 1.305908013786085e+17, 1.305908013907964e+17, 1.305908014029842e+17, 1.30590801415172e+17, 1.30590801427516e+17, 1.305908014397039e+17, 1.305908014518918e+17, 1.305908014640796e+17, 1.305908014762674e+17, 1.305908014884552e+17, 1.305908015006429e+17, 1.305908015129871e+17, 1.305908015251749e+17, 1.305908015373628e+17, 1.305908015497068e+17, 1.305908015618947e+17, 1.305908015740824e+17, 1.305908015862703e+17, 1.305908015986144e+17, 1.305908016108022e+17, 1.305908016229901e+17, 1.305908016351779e+17, 1.30590801647522e+17, 1.305908016597098e+17, 1.305908016718976e+17, 1.305908016840854e+17, 1.305908016962732e+17, 1.305908017086173e+17, 1.305908017208051e+17, 1.30590801732993e+17, 1.305908017451808e+17, 1.305908017573686e+17, 1.305908017695565e+17, 1.305908017817443e+17, 1.305908017940883e+17, 1.305908018062761e+17, 1.30590801818464e+17, 1.305908018308081e+17, 1.305908018429958e+17, 1.305908018551837e+17, 1.305908018673715e+17, 1.305908018797157e+17, 1.305908018919035e+17, 1.305908019040913e+17, 1.305908019162792e+17, 1.305908019284669e+17, 1.30590801940811e+17, 1.305908019529988e+17, 1.305908019651867e+17, 1.305908019773745e+17, 1.305908019895622e+17, 1.305908020017501e+17, 1.305908020139379e+17, 1.305908020262821e+17, 1.305908020384698e+17, 1.305908020506577e+17, 1.305908020628454e+17, 1.305908020751896e+17, 1.305908020873774e+17, 1.305908020995652e+17, 1.305908021117531e+17, 1.305908021239409e+17, 1.305908021362851e+17, 1.305908021484728e+17, 1.305908021606606e+17, 1.305908021728485e+17, 1.305908021851924e+17, 1.305908021973805e+17, 1.30590802209412e+17, 1.305908022217559e+17, 1.305908022339438e+17, 1.305908022461316e+17, 1.305908022583195e+17, 1.305908022706636e+17, 1.305908022826952e+17, 1.305908022950392e+17, 1.30590802307227e+17, 1.305908023194149e+17, 1.305908023317588e+17, 1.305908023439468e+17, 1.305908023561345e+17, 1.305908023683223e+17, 1.305908023805102e+17, 1.305908023928543e+17, 1.305908024050422e+17, 1.3059080241723e+17, 1.305908024294177e+17, 1.305908024416056e+17, 1.305908024537934e+17, 1.305908024661376e+17, 1.305908024783252e+17, 1.305908024905132e+17, 1.305908025027011e+17, 1.305908025148888e+17, 1.305908025270767e+17, 1.305908025394207e+17, 1.305908025516086e+17, 1.305908025637964e+17, 1.305908025759841e+17, 1.30590802588172e+17, 1.30590802600516e+17, 1.305908026127039e+17, 1.305908026248916e+17, 1.305908026370796e+17, 1.305908026494236e+17, 1.305908026616114e+17, 1.305908026739555e+17, 1.305908026861434e+17, 1.305908026983313e+17, 1.30590802710519e+17, 1.305908027227068e+17, 1.305908027348947e+17, 1.305908027472388e+17, 1.305908027594266e+17, 1.305908027716143e+17, 1.305908027838022e+17, 1.305908027961462e+17, 1.305908028083341e+17, 1.30590802820522e+17, 1.305908028327098e+17, 1.305908028448975e+17, 1.305908028570853e+17, 1.305908028692732e+17, 1.305908028814611e+17, 1.305908028938052e+17, 1.30590802905993e+17, 1.305908029181807e+17, 1.305908029303686e+17, 1.305908029425564e+17, 1.305908029547442e+17, 1.305908029670884e+17, 1.305908029792762e+17, 1.305908029914641e+17, 1.30590803003808e+17, 1.305908030159959e+17, 1.305908030281837e+17, 1.305908030405277e+17, 1.305908030527155e+17, 1.305908030649034e+17, 1.305908030770913e+17, 1.305908030892791e+17, 1.305908031016232e+17, 1.305908031138109e+17, 1.305908031259988e+17, 1.305908031383429e+17, 1.305908031505307e+17, 1.305908031627186e+17, 1.305908031749064e+17, 1.305908031872506e+17, 1.305908031994383e+17, 1.305908032116261e+17, 1.305908032238139e+17, 1.305908032360017e+17, 1.305908032481896e+17, 1.305908032603775e+17, 1.305908032727215e+17, 1.305908032849093e+17, 1.305908032970971e+17, 1.30590803309285e+17, 1.305908033214728e+17, 1.305908033336607e+17, 1.305908033460046e+17, 1.305908033581925e+17, 1.305908033703803e+17, 1.305908033825681e+17, 1.30590803394756e+17, 1.305908034069437e+17, 1.305908034191316e+17, 1.305908034313194e+17, 1.305908034435072e+17, 1.305908034556951e+17, 1.305908034678829e+17, 1.305908034800707e+17, 1.305908034922586e+17, 1.305908035046026e+17, 1.305908035167905e+17, 1.305908035289783e+17, 1.305908035413224e+17, 1.30590803553354e+17, 1.305908035655418e+17, 1.30590803577886e+17, 1.305908035900737e+17, 1.305908036022615e+17, 1.305908036146056e+17, 1.305908036267935e+17, 1.305908036389812e+17, 1.30590803651169e+17, 1.305908036635131e+17, 1.305908036757009e+17, 1.305908036878888e+17, 1.305908037000767e+17, 1.305908037122643e+17, 1.305908037244522e+17, 1.3059080373664e+17, 1.305908037489842e+17, 1.30590803761172e+17, 1.305908037733597e+17, 1.305908037855476e+17, 1.305908037977354e+17, 1.305908038099233e+17, 1.305908038222674e+17, 1.305908038344552e+17, 1.305908038466431e+17, 1.305908038588308e+17, 1.305908038710188e+17, 1.305908038833627e+17, 1.305908038955506e+17, 1.305908039077384e+17, 1.305908039199261e+17, 1.305908039322703e+17, 1.305908039444581e+17, 1.30590803956646e+17, 1.305908039688337e+17, 1.305908039811779e+17, 1.305908039933656e+17, 1.305908040055534e+17, 1.305908040177413e+17, 1.305908040300854e+17, 1.305908040422733e+17, 1.305908040544611e+17, 1.305908040666488e+17, 1.305908040788367e+17, 1.305908040911808e+17, 1.305908041033686e+17, 1.305908041155565e+17, 1.305908041277443e+17, 1.305908041399322e+17, 1.305908041522762e+17, 1.30590804164464e+17, 1.305908041766518e+17, 1.305908041889958e+17, 1.305908042011836e+17, 1.305908042133715e+17, 1.305908042255593e+17, 1.305908042377472e+17, 1.305908042500913e+17, 1.30590804262279e+17, 1.305908042744669e+17, 1.305908042866547e+17, 1.305908042988426e+17, 1.305908043110304e+17, 1.305908043232182e+17, 1.305908043354061e+17, 1.3059080434775e+17, 1.30590804359938e+17, 1.305908043721258e+17, 1.305908043843136e+17, 1.305908043965015e+17, 1.305908044088454e+17, 1.305908044210333e+17, 1.305908044332211e+17, 1.305908044454089e+17, 1.30590804457753e+17, 1.305908044699409e+17, 1.305908044821286e+17, 1.305908044944727e+17, 1.305908045065043e+17, 1.305908045188484e+17, 1.305908045310363e+17, 1.305908045432241e+17, 1.305908045554118e+17, 1.305908045675997e+17, 1.305908045797875e+17, 1.305908045919753e+17, 1.305908046043194e+17, 1.305908046165073e+17, 1.305908046286952e+17, 1.305908046410391e+17, 1.30590804653227e+17, 1.305908046654148e+17, 1.305908046776027e+17, 1.305908046897905e+17, 1.305908047021345e+17, 1.305908047143224e+17, 1.305908047265101e+17, 1.305908047386981e+17, 1.305908047508859e+17, 1.3059080476323e+17, 1.305908047754177e+17, 1.305908047876055e+17, 1.305908047997934e+17, 1.305908048119812e+17, 1.305908048243254e+17, 1.305908048365132e+17, 1.305908048487009e+17, 1.305908048610451e+17, 1.305908048732328e+17, 1.305908048854207e+17, 1.305908048976084e+17, 1.305908049097964e+17, 1.305908049221404e+17, 1.305908049343282e+17, 1.305908049465161e+17, 1.305908049587039e+17, 1.305908049708916e+17, 1.305908049830796e+17, 1.305908049954236e+17, 1.305908050076114e+17, 1.305908050197992e+17, 1.305908050319871e+17, 1.305908050441748e+17, 1.305908050563628e+17, 1.305908050687068e+17, 1.305908050808946e+17, 1.305908050930825e+17, 1.305908051052703e+17, 1.305908051174582e+17, 1.305908051298022e+17, 1.3059080514199e+17, 1.305908051541778e+17, 1.305908051663657e+17, 1.305908051785536e+17, 1.305908051908975e+17, 1.305908052030854e+17, 1.305908052152732e+17, 1.305908052276174e+17, 1.305908052398052e+17, 1.30590805251993e+17, 1.305908052641807e+17, 1.305908052763685e+17, 1.305908052887127e+17, 1.305908053009005e+17, 1.305908053130884e+17, 1.305908053252762e+17, 1.305908053374639e+17, 1.305908053496518e+17, 1.305908053618396e+17, 1.305908053741838e+17, 1.305908053863716e+17, 1.305908053985592e+17, 1.305908054107473e+17, 1.30590805422935e+17, 1.305908054352791e+17, 1.305908054474669e+17, 1.305908054596547e+17, 1.305908054718426e+17, 1.305908054840303e+17, 1.305908054962182e+17, 1.305908055085623e+17, 1.305908055207501e+17, 1.30590805532938e+17, 1.305908055451258e+17, 1.305908055573137e+17, 1.305908055695014e+17, 1.305908055818455e+17, 1.305908055940333e+17, 1.305908056062211e+17, 1.30590805618409e+17, 1.30590805630753e+17, 1.305908056429409e+17, 1.305908056551287e+17, 1.305908056673165e+17, 1.305908056796605e+17, 1.305908056918484e+17, 1.305908057040362e+17, 1.30590805716224e+17, 1.305908057284119e+17, 1.30590805740756e+17, 1.305908057529439e+17, 1.305908057651316e+17, 1.305908057773194e+17, 1.305908057895073e+17, 1.305908058018513e+17, 1.305908058140392e+17, 1.305908058262269e+17, 1.305908058384147e+17, 1.305908058506026e+17, 1.305908058627904e+17, 1.305908058751346e+17, 1.305908058873224e+17, 1.305908058995101e+17, 1.30590805911698e+17, 1.305908059238858e+17, 1.305908059360737e+17, 1.305908059484177e+17, 1.305908059606056e+17, 1.305908059727935e+17, 1.305908059849812e+17, 1.30590805997169e+17, 1.305908060095131e+17, 1.30590806021701e+17, 1.305908060338888e+17, 1.30590806046233e+17, 1.305908060584206e+17, 1.305908060706085e+17, 1.305908060827963e+17, 1.305908060949842e+17, 1.30590806107172e+17, 1.30590806119516e+17, 1.305908061317039e+17, 1.305908061438917e+17, 1.305908061560795e+17, 1.305908061682674e+17, 1.305908061804552e+17, 1.305908061926429e+17, 1.30590806204987e+17, 1.305908062171749e+17, 1.305908062293628e+17, 1.305908062415506e+17, 1.305908062537384e+17, 1.305908062660824e+17, 1.305908062782702e+17, 1.305908062904581e+17, 1.305908063026459e+17, 1.305908063148338e+17, 1.305908063271777e+17, 1.305908063393656e+17, 1.305908063515535e+17, 1.305908063637412e+17, 1.305908063759291e+17, 1.305908063881169e+17, 1.305908064004611e+17, 1.305908064126488e+17, 1.305908064248366e+17, 1.305908064371808e+17, 1.305908064492123e+17, 1.305908064615565e+17, 1.305908064737443e+17, 1.30590806485932e+17, 1.305908064981199e+17, 1.305908065103077e+17, 1.305908065224956e+17, 1.305908065346834e+17, 1.305908065470275e+17, 1.305908065592152e+17, 1.30590806571403e+17, 1.305908065837472e+17, 1.30590806595935e+17, 1.305908066081229e+17, 1.305908066203107e+17, 1.305908066324984e+17, 1.305908066448425e+17, 1.305908066570304e+17, 1.305908066692182e+17, 1.30590806681406e+17, 1.305908066935939e+17, 1.305908067057816e+17, 1.305908067181258e+17, 1.305908067303136e+17, 1.305908067425014e+17, 1.305908067546893e+17, 1.305908067668771e+17, 1.305908067792212e+17, 1.30590806791409e+17, 1.305908068035967e+17, 1.305908068157846e+17, 1.305908068281286e+17, 1.305908068403165e+17, 1.305908068525043e+17, 1.305908068646921e+17, 1.3059080687688e+17, 1.305908068892241e+17, 1.30590806901412e+17, 1.305908069135997e+17, 1.305908069257875e+17, 1.305908069379753e+17, 1.305908069503195e+17, 1.305908069625073e+17, 1.30590806974695e+17, 1.305908069868829e+17, 1.30590806999227e+17, 1.305908070114149e+17, 1.305908070236027e+17, 1.305908070357905e+17, 1.305908070479784e+17, 1.305908070601661e+17, 1.305908070723539e+17, 1.30590807084698e+17, 1.305908070968859e+17, 1.305908071090737e+17, 1.305908071212614e+17, 1.305908071334493e+17, 1.305908071456371e+17, 1.305908071578249e+17, 1.305908071701691e+17, 1.305908071823567e+17, 1.305908071945446e+17, 1.305908072067325e+17, 1.305908072189203e+17, 1.305908072311081e+17, 1.305908072434522e+17, 1.305908072556401e+17, 1.305908072678278e+17, 1.305908072800157e+17, 1.305908072922035e+17, 1.305908073045476e+17, 1.305908073167355e+17, 1.305908073290796e+17, 1.305908073411112e+17, 1.305908073532989e+17, 1.30590807365643e+17, 1.305908073778308e+17, 1.305908073900187e+17, 1.305908074022066e+17, 1.305908074143944e+17, 1.305908074265821e+17, 1.305908074389262e+17, 1.30590807451114e+17, 1.305908074633019e+17, 1.305908074754897e+17, 1.305908074876776e+17, 1.305908074998653e+17, 1.305908075122094e+17, 1.305908075243972e+17, 1.30590807536585e+17, 1.305908075489292e+17, 1.305908075611169e+17, 1.305908075733048e+17, 1.305908075854926e+17, 1.305908075976804e+17, 1.305908076100244e+17, 1.305908076222122e+17, 1.305908076344003e+17, 1.30590807646588e+17, 1.305908076587758e+17, 1.305908076709636e+17, 1.305908076833076e+17, 1.305908076954956e+17, 1.305908077076833e+17, 1.305908077198712e+17, 1.305908077322152e+17, 1.305908077444031e+17, 1.30590807756591e+17, 1.305908077687786e+17, 1.305908077809665e+17, 1.305908077933106e+17, 1.305908078053422e+17, 1.305908078176863e+17, 1.30590807829874e+17, 1.30590807842062e+17, 1.30590807854406e+17, 1.305908078665938e+17, 1.305908078787817e+17, 1.305908078909695e+17, 1.305908079031574e+17, 1.305908079153452e+17, 1.305908079275331e+17, 1.305908079397208e+17, 1.305908079519086e+17, 1.305908079640965e+17, 1.305908079762843e+17, 1.305908079886284e+17, 1.305908080008161e+17, 1.30590808013004e+17, 1.305908080251918e+17, 1.305908080373796e+17, 1.305908080495675e+17, 1.305908080619116e+17, 1.305908080740995e+17, 1.305908080862872e+17, 1.305908080984749e+17, 1.305908081106628e+17, 1.305908081228507e+17, 1.305908081350385e+17, 1.305908081472264e+17, 1.305908081594141e+17, 1.305908081717582e+17, 1.30590808183946e+17, 1.305908081961339e+17, 1.305908082083217e+17, 1.305908082205094e+17, 1.305908082326973e+17, 1.305908082450414e+17, 1.305908082572293e+17, 1.305908082694171e+17, 1.305908082816049e+17, 1.305908082937928e+17, 1.305908083059805e+17, 1.305908083181683e+17, 1.305908083305124e+17, 1.305908083427003e+17, 1.305908083548881e+17, 1.305908083670758e+17, 1.3059080837942e+17, 1.305908083916077e+17, 1.305908084037957e+17, 1.305908084159835e+17, 1.305908084281713e+17, 1.305908084403592e+17, 1.305908084525468e+17, 1.30590808464891e+17, 1.305908084770788e+17, 1.305908084892667e+17, 1.305908085014545e+17, 1.305908085136422e+17, 1.305908085258301e+17, 1.305908085381742e+17, 1.305908085503621e+17, 1.305908085625499e+17, 1.305908085747377e+17, 1.305908085869256e+17, 1.305908085991133e+17, 1.305908086114574e+17, 1.305908086236452e+17, 1.305908086359892e+17, 1.30590808648177e+17, 1.305908086602086e+17, 1.305908086723965e+17, 1.305908086847406e+17, 1.305908086969284e+17, 1.305908087091162e+17, 1.305908087213039e+17, 1.305908087334918e+17, 1.305908087456797e+17, 1.305908087578675e+17, 1.305908087702116e+17, 1.305908087823994e+17, 1.305908087945873e+17, 1.30590808806775e+17, 1.305908088189629e+17, 1.30590808831307e+17, 1.305908088434948e+17, 1.305908088556826e+17, 1.305908088680268e+17, 1.305908088802145e+17, 1.305908088922461e+17, 1.305908089044339e+17, 1.30590808916778e+17, 1.305908089289658e+17, 1.305908089413098e+17, 1.305908089534977e+17, 1.305908089656855e+17, 1.305908089778733e+17, 1.305908089900612e+17, 1.305908090024052e+17, 1.30590809014593e+17, 1.305908090267809e+17, 1.305908090389687e+17, 1.305908090511566e+17, 1.305908090635005e+17, 1.305908090756884e+17, 1.305908090878764e+17, 1.305908091002204e+17, 1.305908091122519e+17, 1.305908091244397e+17, 1.305908091367839e+17, 1.305908091489716e+17, 1.305908091611594e+17, 1.305908091733473e+17, 1.305908091856914e+17, 1.305908091978792e+17, 1.305908092100669e+17, 1.305908092222548e+17, 1.305908092345989e+17, 1.305908092467868e+17, 1.305908092589746e+17, 1.305908092711624e+17, 1.305908092833503e+17, 1.305908092956943e+17, 1.305908093078822e+17, 1.305908093200699e+17, 1.305908093322578e+17, 1.305908093444456e+17, 1.305908093566335e+17, 1.305908093689775e+17, 1.305908093811653e+17, 1.305908093933532e+17, 1.30590809405541e+17, 1.305908094177288e+17, 1.305908094299167e+17, 1.305908094422606e+17, 1.305908094544485e+17, 1.305908094666363e+17, 1.305908094788241e+17, 1.30590809491012e+17, 1.30590809503356e+17, 1.305908095155439e+17, 1.305908095277317e+17, 1.305908095399195e+17, 1.305908095521074e+17, 1.305908095642952e+17, 1.305908095764831e+17, 1.30590809588827e+17, 1.305908096010149e+17, 1.305908096132027e+17, 1.305908096253906e+17, 1.305908096375785e+17, 1.305908096497661e+17, 1.305908096621102e+17, 1.30590809674298e+17, 1.305908096864859e+17, 1.305908096986738e+17, 1.305908097108616e+17, 1.305908097232056e+17, 1.305908097353934e+17, 1.305908097475813e+17, 1.305908097599254e+17, 1.305908097721133e+17, 1.305908097843011e+17, 1.305908097964888e+17, 1.305908098086767e+17, 1.305908098210207e+17, 1.305908098332086e+17, 1.305908098453965e+17, 1.305908098575841e+17, 1.30590809869772e+17, 1.305908098819598e+17, 1.30590809894304e+17, 1.305908099064918e+17, 1.305908099186796e+17, 1.305908099308673e+17, 1.305908099430551e+17, 1.30590809955243e+17, 1.305908099675871e+17, 1.30590809979775e+17, 1.305908099919628e+17, 1.305908100041505e+17, 1.305908100163384e+17, 1.305908100286825e+17, 1.305908100408704e+17, 1.305908100530582e+17, 1.305908100654022e+17, 1.3059081007759e+17, 1.305908100897779e+17, 1.305908101019657e+17, 1.305908101143098e+17, 1.305908101264975e+17, 1.305908101386853e+17, 1.305908101508732e+17, 1.305908101630611e+17, 1.305908101754052e+17, 1.30590810187593e+17, 1.305908101997807e+17, 1.305908102119686e+17, 1.305908102241564e+17, 1.305908102365006e+17, 1.305908102486884e+17, 1.305908102610324e+17, 1.305908102732202e+17, 1.30590810285408e+17, 1.305908102975959e+17, 1.305908103097837e+17, 1.305908103221279e+17, 1.305908103343156e+17, 1.305908103465034e+17, 1.305908103586912e+17, 1.30590810370879e+17, 1.30590810383067e+17, 1.305908103954109e+17, 1.305908104075988e+17, 1.305908104199428e+17, 1.305908104321307e+17, 1.305908104443186e+17, 1.305908104565064e+17, 1.305908104688504e+17, 1.305908104810382e+17, 1.305908104932261e+17, 1.305908105054139e+17, 1.305908105177581e+17, 1.305908105299457e+17, 1.305908105421336e+17, 1.305908105543214e+17, 1.305908105665092e+17, 1.305908105788534e+17, 1.305908105910412e+17, 1.305908106032291e+17, 1.30590810615573e+17, 1.305908106277609e+17, 1.305908106399487e+17, 1.305908106521366e+17, 1.305908106643245e+17, 1.305908106726058e+17, 1.305908106847936e+17, 1.305908106969815e+17, 1.305908107091693e+17, 1.305908107213571e+17, 1.305908107337012e+17, 1.30590810745889e+17, 1.305908107540142e+17, 1.305908107662021e+17, 1.305908107783899e+17, 1.305908107905777e+17, 1.305908108029217e+17, 1.305908108151096e+17, 1.305908108272974e+17, 1.305908108396415e+17, 1.305908108518294e+17, 1.305908108640172e+17, 1.305908108762051e+17, 1.30590810888549e+17, 1.305908109007369e+17, 1.305908109088621e+17, 1.3059081092105e+17, 1.30590810933394e+17, 1.305908109455818e+17, 1.305908109537071e+17, 1.305908109660511e+17, 1.30590810978239e+17, 1.305908109904269e+17, 1.305908110026145e+17, 1.305908110148024e+17, 1.305908110271465e+17, 1.305908110393343e+17, 1.30590811051522e+17, 1.3059081106371e+17, 1.305908110758977e+17, 1.305908110882419e+17, 1.305908111004297e+17, 1.305908111126175e+17, 1.305908111249617e+17, 1.305908111371494e+17, 1.305908111493373e+17, 1.305908111615251e+17, 1.305908111738692e+17, 1.30590811186057e+17, 1.305908111982447e+17, 1.305908112104326e+17, 1.305908112226204e+17, 1.305908112348083e+17, 1.305908112471523e+17, 1.305908112593402e+17, 1.305908112715279e+17, 1.305908112837157e+17, 1.305908112959036e+17, 1.305908113080914e+17, 1.305908113204356e+17, 1.305908113326234e+17, 1.305908113448111e+17, 1.30590811356999e+17, 1.305908113691868e+17, 1.305908113813747e+17, 1.305908113935625e+17, 1.305908114059066e+17, 1.305908114180945e+17, 1.305908114302821e+17, 1.305908114423137e+17, 1.305908114546579e+17, 1.305908114668457e+17, 1.305908114790336e+17, 1.305908114913775e+17, 1.305908115035654e+17, 1.305908115155969e+17, 1.30590811527941e+17, 1.305908115401289e+17, 1.305908115523167e+17, 1.305908115646607e+17, 1.305908115768485e+17, 1.305908115890364e+17, 1.305908116012242e+17, 1.30590811613412e+17, 1.305908116255999e+17, 1.305908116377876e+17, 1.305908116501318e+17, 1.305908116623196e+17, 1.305908116745074e+17, 1.305908116866953e+17, 1.305908116990394e+17, 1.305908117112271e+17, 1.30590811723415e+17, 1.305908117356028e+17, 1.305908117477907e+17, 1.305908117599784e+17, 1.305908117723226e+17, 1.305908117845103e+17, 1.305908117966982e+17, 1.30590811808886e+17, 1.305908118210738e+17, 1.305908118332616e+17, 1.305908118456056e+17, 1.305908118577935e+17, 1.305908118699813e+17, 1.305908118823255e+17, 1.305908118945133e+17, 1.305908119067011e+17, 1.30590811918889e+17, 1.30590811931233e+17, 1.305908119434208e+17, 1.305908119556086e+17, 1.305908119677965e+17, 1.305908119799843e+17, 1.305908119923284e+17, 1.305908120045162e+17, 1.30590812016704e+17, 1.305908120288919e+17, 1.305908120410797e+17, 1.305908120532675e+17, 1.305908120656115e+17, 1.305908120777994e+17, 1.305908120899872e+17, 1.30590812102175e+17, 1.305908121143629e+17, 1.305908121267069e+17, 1.305908121388948e+17, 1.305908121510826e+17, 1.305908121632704e+17, 1.305908121754583e+17, 1.305908121876461e+17, 1.305908121998339e+17, 1.305908122121779e+17, 1.305908122243657e+17, 1.305908122365536e+17, 1.305908122487414e+17, 1.305908122609293e+17, 1.305908122731172e+17, 1.305908122854611e+17, 1.30590812297649e+17, 1.305908123098367e+17, 1.305908123220246e+17, 1.305908123343686e+17, 1.305908123465565e+17, 1.305908123587443e+17, 1.305908123710885e+17, 1.305908123832762e+17, 1.305908123954641e+17, 1.30590812407652e+17, 1.305908124198397e+17, 1.305908124320275e+17, 1.305908124443716e+17, 1.305908124565595e+17, 1.305908124687473e+17, 1.30590812480935e+17, 1.305908124931229e+17, 1.305908125053107e+17, 1.305908125176548e+17, 1.305908125298426e+17, 1.305908125420305e+17, 1.305908125542184e+17, 1.305908125664061e+17, 1.305908125787502e+17, 1.30590812590938e+17, 1.305908126031259e+17, 1.305908126153137e+17, 1.305908126276577e+17, 1.305908126398456e+17, 1.305908126520334e+17, 1.305908126642213e+17, 1.305908126764091e+17, 1.305908126887532e+17, 1.305908127009409e+17, 1.305908127131287e+17, 1.305908127253166e+17, 1.305908127376605e+17, 1.305908127498486e+17, 1.305908127620364e+17, 1.305908127742241e+17, 1.305908127864119e+17, 1.30590812798756e+17, 1.305908128109439e+17, 1.305908128231316e+17, 1.305908128353196e+17, 1.305908128475073e+17, 1.305908128596951e+17, 1.30590812871883e+17, 1.305908128842271e+17, 1.30590812896415e+17, 1.305908129086028e+17, 1.305908129207905e+17, 1.305908129329783e+17, 1.305908129453224e+17, 1.305908129575103e+17, 1.30590812969698e+17, 1.305908129820421e+17, 1.305908129942299e+17, 1.305908130064178e+17, 1.305908130186057e+17, 1.305908130307933e+17, 1.305908130431375e+17, 1.305908130553253e+17, 1.305908130675132e+17, 1.30590813079701e+17, 1.305908130918888e+17, 1.305908131040767e+17, 1.305908131164207e+17, 1.305908131286085e+17, 1.305908131407964e+17, 1.305908131529842e+17, 1.305908131651721e+17, 1.305908131773599e+17, 1.305908131897039e+17, 1.305908132018917e+17, 1.305908132140796e+17, 1.305908132262674e+17, 1.305908132384552e+17, 1.305908132506431e+17, 1.30590813262987e+17, 1.305908132751749e+17, 1.305908132873627e+17, 1.305908132995506e+17, 1.305908133117384e+17, 1.305908133239261e+17, 1.305908133362703e+17, 1.305908133484581e+17, 1.30590813360646e+17, 1.305908133728338e+17, 1.305908133850216e+17, 1.305908133973656e+17, 1.305908134095534e+17, 1.305908134217414e+17, 1.305908134339292e+17, 1.30590813446117e+17, 1.305908134583048e+17, 1.305908134704925e+17, 1.305908134828367e+17, 1.305908134950245e+17, 1.305908135073686e+17, 1.305908135195564e+17, 1.305908135317443e+17, 1.30590813543932e+17, 1.305908135561198e+17, 1.30590813568464e+17, 1.305908135806518e+17, 1.305908135928397e+17, 1.305908136050275e+17, 1.305908136173715e+17, 1.305908136295594e+17, 1.305908136417472e+17, 1.30590813653935e+17, 1.305908136661228e+17, 1.305908136784669e+17, 1.305908136906547e+17, 1.305908137028425e+17, 1.305908137150304e+17, 1.305908137273745e+17, 1.305908137395622e+17, 1.3059081375175e+17, 1.305908137639379e+17, 1.305908137761257e+17, 1.305908137883135e+17, 1.305908138006577e+17, 1.305908138128454e+17, 1.305908138250333e+17, 1.305908138372211e+17, 1.305908138494089e+17, 1.30590813861753e+17, 1.305908138737846e+17, 1.305908138861288e+17, 1.305908138983164e+17, 1.305908139105043e+17, 1.305908139226921e+17, 1.305908139350362e+17, 1.305908139472239e+17, 1.305908139594118e+17, 1.305908139715997e+17, 1.305908139837874e+17, 1.305908139959753e+17, 1.305908140081632e+17, 1.305908140205071e+17, 1.30590814032695e+17, 1.305908140448828e+17, 1.305908140570707e+17, 1.305908140692585e+17, 1.305908140814463e+17, 1.305908140936342e+17, 1.30590814105822e+17, 1.305908141180097e+17, 1.305908141301976e+17, 1.305908141425417e+17, 1.305908141547296e+17, 1.305908141669174e+17, 1.305908141792614e+17, 1.305908141912931e+17, 1.305908142034808e+17, 1.305908142156687e+17, 1.305908142280128e+17, 1.305908142402006e+17, 1.305908142525446e+17, 1.305908142647324e+17, 1.305908142769202e+17, 1.30590814289108e+17, 1.30590814301296e+17, 1.305908143134838e+17, 1.305908143258278e+17, 1.305908143378593e+17, 1.305908143500471e+17, 1.305908143623913e+17, 1.305908143745791e+17, 1.30590814386767e+17, 1.30590814399111e+17, 1.305908144112988e+17, 1.305908144234867e+17, 1.305908144356745e+17, 1.305908144480186e+17, 1.305908144602063e+17, 1.305908144725504e+17, 1.305908144847382e+17, 1.305908144969262e+17, 1.30590814509114e+17, 1.305908145213018e+17, 1.305908145334895e+17, 1.305908145456773e+17, 1.305908145580215e+17, 1.305908145702093e+17, 1.305908145823972e+17, 1.30590814594585e+17, 1.30590814606929e+17, 1.305908146191169e+17, 1.305908146313047e+17, 1.305908146434926e+17, 1.305908146556804e+17, 1.305908146680244e+17, 1.305908146802122e+17, 1.305908146924e+17, 1.305908147045879e+17, 1.305908147167757e+17, 1.305908147289636e+17, 1.305908147413075e+17, 1.305908147534954e+17, 1.305908147656833e+17, 1.305908147778711e+17, 1.305908147900589e+17, 1.305908148024029e+17, 1.305908148145908e+17, 1.305908148267786e+17, 1.305908148389664e+17, 1.305908148513106e+17, 1.305908148634984e+17, 1.305908148756863e+17, 1.30590814887874e+17, 1.305908149002181e+17, 1.305908149124059e+17, 1.305908149245937e+17, 1.305908149367816e+17, 1.305908149489693e+17, 1.305908149611572e+17, 1.305908149735012e+17, 1.305908149856891e+17, 1.305908149978769e+17, 1.305908150100646e+17, 1.305908150222525e+17, 1.305908150345966e+17, 1.305908150467845e+17, 1.305908150589723e+17, 1.305908150713164e+17, 1.305908150835041e+17, 1.30590815095692e+17, 1.305908151078799e+17, 1.305908151202239e+17, 1.305908151324118e+17, 1.305908151445996e+17, 1.305908151567873e+17, 1.305908151689752e+17, 1.305908151813193e+17, 1.305908151935071e+17, 1.305908152056948e+17, 1.30590815218039e+17, 1.305908152302268e+17, 1.305908152424147e+17, 1.305908152547588e+17, 1.305908152669466e+17, 1.305908152791343e+17, 1.305908152913221e+17, 1.305908153035101e+17, 1.305908153156979e+17, 1.305908153278857e+17, 1.305908153402298e+17, 1.305908153524175e+17, 1.305908153646054e+17, 1.305908153767932e+17, 1.305908153889811e+17, 1.305908154011689e+17, 1.30590815413513e+17, 1.305908154257007e+17, 1.305908154378885e+17, 1.305908154500764e+17, 1.305908154622642e+17, 1.305908154746084e+17, 1.305908154867962e+17, 1.305908154989839e+17, 1.305908155111718e+17, 1.305908155233596e+17, 1.305908155355475e+17, 1.305908155478915e+17, 1.305908155600794e+17, 1.305908155722673e+17, 1.30590815584455e+17, 1.305908155966428e+17, 1.305908156088306e+17, 1.305908156211747e+17, 1.305908156333626e+17, 1.305908156455503e+17, 1.305908156577382e+17, 1.30590815669926e+17, 1.305908156821138e+17, 1.305908156944579e+17, 1.305908157066458e+17, 1.305908157188335e+17, 1.305908157310213e+17, 1.305908157432092e+17, 1.305908157555533e+17, 1.305908157677412e+17, 1.30590815779929e+17, 1.305908157921167e+17, 1.305908158044608e+17, 1.305908158166486e+17, 1.305908158288365e+17, 1.305908158410244e+17, 1.305908158532122e+17, 1.305908158655562e+17, 1.30590815877744e+17, 1.305908158899318e+17, 1.305908159021197e+17, 1.305908159143076e+17, 1.305908159266515e+17, 1.305908159388394e+17, 1.305908159510272e+17, 1.30590815963215e+17, 1.305908159754029e+17, 1.305908159877469e+17, 1.305908159999348e+17, 1.305908160121226e+17, 1.305908160243104e+17, 1.305908160364983e+17, 1.305908160488422e+17, 1.305908160610301e+17, 1.305908160732179e+17, 1.30590816085562e+17, 1.305908160977499e+17, 1.305908161099377e+17, 1.305908161221256e+17, 1.305908161344696e+17, 1.305908161466574e+17, 1.305908161588452e+17, 1.305908161710331e+17, 1.305908161832209e+17, 1.305908161954086e+17, 1.305908162077528e+17, 1.305908162199406e+17, 1.305908162321285e+17, 1.305908162443163e+17, 1.305908162565041e+17, 1.30590816268692e+17, 1.30590816281036e+17, 1.305908162932238e+17, 1.305908163054117e+17, 1.305908163175995e+17, 1.305908163297873e+17, 1.30590816341975e+17, 1.305908163543191e+17, 1.305908163665069e+17, 1.305908163786949e+17, 1.305908163908827e+17, 1.305908164030705e+17, 1.305908164152582e+17, 1.30590816427446e+17, 1.305908164397902e+17, 1.30590816451978e+17, 1.305908164641659e+17, 1.3059081647651e+17, 1.305908164885414e+17, 1.305908165008856e+17, 1.305908165130734e+17, 1.305908165252613e+17, 1.305908165374491e+17, 1.305908165496369e+17, 1.305908165619809e+17, 1.305908165741687e+17, 1.305908165863566e+17, 1.305908165985444e+17, 1.305908166107323e+17, 1.305908166230762e+17, 1.305908166352641e+17, 1.30590816647452e+17, 1.305908166596398e+17, 1.305908166718277e+17, 1.305908166840154e+17, 1.305908166963596e+17, 1.305908167085473e+17, 1.305908167207351e+17, 1.30590816732923e+17, 1.305908167452671e+17, 1.30590816757455e+17, 1.305908167696428e+17, 1.305908167818305e+17, 1.305908167940184e+17, 1.305908168062062e+17, 1.305908168185503e+17, 1.30590816830738e+17, 1.30590816842926e+17, 1.305908168551137e+17, 1.305908168673015e+17, 1.305908168794894e+17, 1.305908168918333e+17, 1.305908169040214e+17, 1.305908169162092e+17, 1.305908169283969e+17, 1.30590816940741e+17, 1.305908169527725e+17, 1.305908169651167e+17, 1.305908169773044e+17, 1.305908169894924e+17, 1.305908170016801e+17, 1.305908170140242e+17, 1.30590817026212e+17, 1.305908170383999e+17, 1.305908170507439e+17, 1.305908170629317e+17, 1.305908170751196e+17, 1.305908170873074e+17, 1.305908170994952e+17, 1.305908171118392e+17, 1.305908171240271e+17, 1.305908171362149e+17, 1.305908171484027e+17, 1.305908171605906e+17, 1.305908171727785e+17, 1.305908171851226e+17, 1.305908171973103e+17, 1.305908172094981e+17, 1.30590817221686e+17, 1.3059081723403e+17, 1.30590817246218e+17, 1.305908172584058e+17, 1.305908172705935e+17, 1.305908172827814e+17, 1.305908172951254e+17, 1.305908173073133e+17, 1.305908173195011e+17, 1.305908173318451e+17, 1.305908173440329e+17, 1.305908173562208e+17, 1.305908173684086e+17, 1.305908173805965e+17, 1.305908173927843e+17, 1.305908174051283e+17, 1.305908174173162e+17, 1.30590817429504e+17, 1.305908174416918e+17, 1.305908174538797e+17, 1.305908174662237e+17, 1.305908174784115e+17, 1.305908174905993e+17, 1.305908175027872e+17, 1.305908175149751e+17, 1.30590817527319e+17, 1.305908175395069e+17, 1.305908175516947e+17, 1.305908175638825e+17, 1.305908175762266e+17, 1.305908175884145e+17, 1.305908176006022e+17, 1.305908176129464e+17, 1.305908176251342e+17, 1.30590817637322e+17, 1.305908176496662e+17, 1.30590817661854e+17, 1.305908176740417e+17, 1.305908176862295e+17, 1.305908176984173e+17, 1.305908177106053e+17, 1.305908177227931e+17, 1.305908177351372e+17, 1.305908177473249e+17, 1.305908177595127e+17, 1.305908177718568e+17, 1.305908177840447e+17, 1.305908177962324e+17, 1.305908178084202e+17, 1.305908178206081e+17, 1.305908178329522e+17, 1.305908178451401e+17, 1.305908178573279e+17, 1.305908178695156e+17, 1.305908178817036e+17, 1.305908178938913e+17, 1.305908179062354e+17, 1.305908179184233e+17, 1.305908179306111e+17, 1.305908179427988e+17, 1.305908179549866e+17, 1.305908179673308e+17, 1.305908179795186e+17, 1.305908179917065e+17, 1.305908180038943e+17, 1.305908180160819e+17, 1.305908180282698e+17, 1.305908180404577e+17, 1.305908180528018e+17, 1.305908180649896e+17, 1.305908180771773e+17, 1.305908180893652e+17, 1.30590818101553e+17, 1.305908181138972e+17, 1.30590818126085e+17, 1.305908181382728e+17, 1.305908181504607e+17, 1.305908181628047e+17, 1.305908181749926e+17, 1.305908181871804e+17, 1.305908181993682e+17, 1.30590818211556e+17, 1.305908182239002e+17, 1.305908182360878e+17, 1.305908182482757e+17, 1.305908182604636e+17, 1.305908182728076e+17, 1.305908182849955e+17, 1.305908182971832e+17, 1.305908183093711e+17, 1.305908183215589e+17, 1.305908183337467e+17, 1.305908183460909e+17, 1.305908183582787e+17, 1.305908183704666e+17, 1.305908183826543e+17, 1.305908183948421e+17, 1.305908184071862e+17, 1.30590818419374e+17, 1.305908184315619e+17, 1.305908184437496e+17, 1.305908184559374e+17, 1.305908184681253e+17, 1.305908184804694e+17, 1.305908184926572e+17, 1.305908185048449e+17, 1.305908185170328e+17, 1.305908185292207e+17, 1.305908185415648e+17, 1.305908185537526e+17, 1.305908185659404e+17, 1.305908185781283e+17, 1.305908185904723e+17, 1.305908186026602e+17, 1.30590818614848e+17, 1.305908186270358e+17, 1.305908186392237e+17, 1.305908186515676e+17, 1.305908186637555e+17, 1.305908186759433e+17, 1.305908186881312e+17, 1.30590818700319e+17, 1.30590818712663e+17, 1.305908187248509e+17, 1.305908187370387e+17, 1.305908187492266e+17, 1.305908187614143e+17, 1.305908187737585e+17, 1.305908187859462e+17, 1.30590818798134e+17, 1.305908188104782e+17, 1.30590818822666e+17, 1.305908188348539e+17, 1.305908188470417e+17, 1.305908188592294e+17, 1.305908188715735e+17, 1.305908188837613e+17, 1.305908188959492e+17, 1.30590818908137e+17, 1.305908189203249e+17, 1.305908189325126e+17, 1.305908189448567e+17, 1.305908189570445e+17, 1.305908189692323e+17, 1.305908189814202e+17, 1.305908189936079e+17, 1.305908190057958e+17, 1.305908190181399e+17, 1.305908190303277e+17, 1.305908190425156e+17, 1.305908190547034e+17, 1.305908190668913e+17, 1.305908190792352e+17, 1.305908190914231e+17, 1.305908191036109e+17, 1.305908191157987e+17, 1.305908191281427e+17, 1.305908191403306e+17, 1.305908191525184e+17, 1.305908191648625e+17, 1.305908191770504e+17, 1.305908191892381e+17, 1.305908192014259e+17, 1.305908192136138e+17, 1.305908192258016e+17, 1.305908192381457e+17, 1.305908192503334e+17, 1.305908192625213e+17, 1.305908192747091e+17, 1.305908192868969e+17, 1.30590819299241e+17, 1.305908193114289e+17, 1.305908193236166e+17, 1.305908193358044e+17, 1.305908193479923e+17, 1.305908193601801e+17, 1.305908193725243e+17, 1.305908193847121e+17, 1.305908193968998e+17, 1.305908194090876e+17, 1.305908194212755e+17, 1.305908194336196e+17, 1.305908194458074e+17, 1.305908194579953e+17, 1.30590819470183e+17, 1.305908194823707e+17, 1.305908194945586e+17, 1.305908195069027e+17, 1.305908195190906e+17, 1.305908195312783e+17, 1.305908195436225e+17, 1.305908195558103e+17, 1.305908195679981e+17, 1.305908195801859e+17, 1.305908195925299e+17, 1.305908196047177e+17, 1.305908196169055e+17, 1.305908196290935e+17, 1.305908196414374e+17, 1.305908196536253e+17, 1.305908196658131e+17, 1.305908196781573e+17, 1.30590819690345e+17, 1.305908197025329e+17, 1.305908197147206e+17, 1.305908197269085e+17, 1.305908197392526e+17, 1.305908197514404e+17, 1.305908197636283e+17, 1.305908197758161e+17, 1.305908197880037e+17, 1.305908198003479e+17, 1.305908198125357e+17, 1.305908198247236e+17, 1.305908198369114e+17, 1.305908198492556e+17, 1.305908198614433e+17, 1.305908198736311e+17, 1.305908198858189e+17, 1.305908198980067e+17, 1.305908199103507e+17, 1.305908199225386e+17, 1.305908199347265e+17, 1.305908199469143e+17, 1.305908199591021e+17, 1.305908199714461e+17, 1.305908199836339e+17, 1.305908199958218e+17, 1.305908200080096e+17, 1.305908200201975e+17, 1.305908200323853e+17, 1.305908200447293e+17, 1.305908200569171e+17, 1.305908200691049e+17, 1.305908200812928e+17, 1.305908200934806e+17, 1.305908201056684e+17, 1.305908201180124e+17, 1.305908201302003e+17, 1.305908201423881e+17, 1.30590820154576e+17, 1.305908201669201e+17, 1.305908201791078e+17, 1.305908201912957e+17, 1.305908202034834e+17, 1.305908202156713e+17, 1.305908202278591e+17, 1.305908202402031e+17, 1.30590820252391e+17, 1.305908202645788e+17, 1.305908202769229e+17, 1.305908202891107e+17, 1.305908203012986e+17, 1.305908203134863e+17, 1.305908203256741e+17, 1.305908203380183e+17, 1.305908203502061e+17, 1.30590820362394e+17, 1.305908203745818e+17, 1.305908203869258e+17, 1.305908203991136e+17, 1.305908204113014e+17, 1.305908204234892e+17, 1.305908204356771e+17, 1.30590820447865e+17, 1.305908204602089e+17, 1.305908204723968e+17, 1.305908204845846e+17, 1.305908204967724e+17, 1.305908205089603e+17, 1.30590820521148e+17, 1.305908205334922e+17, 1.3059082054568e+17, 1.305908205578678e+17, 1.305908205700557e+17, 1.305908205823997e+17, 1.305908205945875e+17, 1.305908206067753e+17, 1.305908206189631e+17, 1.305908206313071e+17, 1.30590820643495e+17, 1.305908206556828e+17, 1.305908206678706e+17, 1.305908206800585e+17, 1.305908206922463e+17, 1.305908207045903e+17, 1.305908207167781e+17, 1.30590820728966e+17, 1.305908207411539e+17, 1.305908207533417e+17, 1.305908207656858e+17, 1.305908207778735e+17, 1.305908207900613e+17, 1.305908208022491e+17, 1.30590820814437e+17, 1.305908208266248e+17, 1.305908208388127e+17, 1.305908208511567e+17, 1.305908208633445e+17, 1.305908208755324e+17, 1.305908208877202e+17, 1.30590820899908e+17, 1.30590820912252e+17, 1.305908209244399e+17, 1.305908209366278e+17, 1.305908209488155e+17, 1.305908209610034e+17, 1.305908209733473e+17, 1.305908209855352e+17, 1.30590820997723e+17, 1.305908210100672e+17, 1.30590821022255e+17, 1.305908210344428e+17, 1.305908210466307e+17, 1.305908210588184e+17, 1.305908210711625e+17, 1.305908210833503e+17, 1.305908210955382e+17, 1.30590821107726e+17, 1.305908211199137e+17, 1.305908211322579e+17, 1.305908211444457e+17, 1.305908211566336e+17, 1.305908211688212e+17, 1.305908211811654e+17, 1.305908211933532e+17, 1.30590821205541e+17, 1.305908212177289e+17, 1.305908212299167e+17, 1.305908212422609e+17, 1.305908212544486e+17, 1.305908212666364e+17, 1.305908212789804e+17, 1.305908212911683e+17, 1.30590821303356e+17, 1.305908213155438e+17, 1.305908213277317e+17, 1.305908213399195e+17, 1.305908213522637e+17, 1.305908213644515e+17, 1.305908213766392e+17, 1.305908213888271e+17, 1.305908214010149e+17, 1.305908214132028e+17, 1.305908214255468e+17, 1.305908214377347e+17, 1.305908214499224e+17, 1.305908214622665e+17, 1.305908214744543e+17, 1.305908214866422e+17, 1.3059082149883e+17, 1.305908215110177e+17, 1.305908215233619e+17, 1.305908215355497e+17, 1.305908215477376e+17, 1.305908215599254e+17, 1.305908215722694e+17, 1.305908215803946e+17, 1.305908215925824e+17, 1.305908216047702e+17, 1.305908216169581e+17, 1.305908216291459e+17, 1.305908216413336e+17, 1.305908216536778e+17, 1.305908216658656e+17, 1.305908216780535e+17, 1.305908216902413e+17, 1.305908217024291e+17, 1.305908217146168e+17, 1.305908217269609e+17, 1.305908217391488e+17, 1.305908217513366e+17, 1.305908217635245e+17, 1.305908217757123e+17, 1.305908217880563e+17, 1.305908218002441e+17, 1.30590821812432e+17, 1.305908218246198e+17, 1.305908218368076e+17, 1.305908218491517e+17, 1.305908218613395e+17, 1.305908218735273e+17, 1.305908218857151e+17, 1.305908218979028e+17, 1.305908219100908e+17, 1.305908219222785e+17, 1.305908219344664e+17, 1.305908219466543e+17, 1.305908219589983e+17, 1.30590821971186e+17, 1.305908219833738e+17, 1.305908219914991e+17, 1.30590822003687e+17, 1.30590822016031e+17, 1.305908220282189e+17, 1.305908220404068e+17, 1.305908220525944e+17, 1.305908220647823e+17, 1.305908220771264e+17, 1.305908220893142e+17, 1.30590822101502e+17, 1.305908221136899e+17, 1.305908221258776e+17, 1.305908221382218e+17, 1.305908221504096e+17, 1.305908221625974e+17, 1.305908221749414e+17, 1.305908221869731e+17, 1.305908221993171e+17, 1.305908222115049e+17, 1.305908222236927e+17, 1.305908222360369e+17, 1.305908222482246e+17, 1.305908222604124e+17, 1.305908222726002e+17, 1.305908222849444e+17, 1.305908222971322e+17, 1.305908223093201e+17, 1.305908223215078e+17, 1.305908223336956e+17, 1.305908223460397e+17, 1.305908223582275e+17, 1.305908223705715e+17, 1.305908223827594e+17, 1.305908223949472e+17, 1.30590822407135e+17, 1.305908224194792e+17, 1.305908224316669e+17, 1.305908224438548e+17, 1.305908224561988e+17, 1.305908224683867e+17, 1.305908224805745e+17, 1.305908224927622e+17, 1.305908225049501e+17, 1.305908225172941e+17, 1.305908225294821e+17, 1.305908225416699e+17, 1.305908225538577e+17, 1.305908225660454e+17, 1.305908225782332e+17, 1.305908225904211e+17, 1.305908226026089e+17, 1.305908226149531e+17, 1.305908226271409e+17, 1.305908226393286e+17, 1.305908226515165e+17, 1.305908226596417e+17, 1.305908226719857e+17, 1.305908226841736e+17, 1.305908226963613e+17, 1.305908227085492e+17, 1.30590822720737e+17, 1.305908227288623e+17, 1.305908227410501e+17, 1.305908227533942e+17, 1.30590822765582e+17, 1.305908227777699e+17, 1.305908227899576e+17, 1.305908228021454e+17, 1.305908228143333e+17, 1.305908228266772e+17, 1.305908228388652e+17, 1.305908228510529e+17, 1.305908228632407e+17, 1.305908228755849e+17, 1.305908228877727e+17, 1.305908228999604e+17, 1.305908229121484e+17, 1.305908229243361e+17, 1.30590822936524e+17, 1.305908229488681e+17, 1.305908229610559e+17, 1.305908229732436e+17, 1.305908229855877e+17, 1.305908229977755e+17, 1.305908230099634e+17, 1.305908230221512e+17, 1.305908230343391e+17, 1.305908230466831e+17, 1.305908230588709e+17, 1.305908230710587e+17, 1.305908230832465e+17, 1.305908230954344e+17, 1.305908231077784e+17, 1.305908231199663e+17, 1.305908231321541e+17, 1.305908231441856e+17, 1.305908231563735e+17, 1.305908231687174e+17, 1.305908231809053e+17, 1.305908231930931e+17, 1.305908232052809e+17, 1.305908232174689e+17, 1.305908232298129e+17, 1.305908232420008e+17, 1.305908232541885e+17, 1.305908232663763e+17, 1.305908232785642e+17, 1.305908232909083e+17, 1.305908233030962e+17, 1.30590823315284e+17, 1.305908233274717e+17, 1.305908233398158e+17, 1.305908233520036e+17, 1.305908233641914e+17, 1.305908233763791e+17, 1.30590823388567e+17, 1.305908234007548e+17, 1.30590823413099e+17, 1.305908234252868e+17, 1.305908234374746e+17, 1.305908234496625e+17, 1.305908234618502e+17, 1.305908234741943e+17, 1.305908234863821e+17, 1.3059082349857e+17, 1.305908235107579e+17, 1.305908235229455e+17, 1.305908235351334e+17, 1.305908235473212e+17, 1.305908235596653e+17, 1.305908235718531e+17, 1.30590823584041e+17, 1.305908235962287e+17, 1.305908236084165e+17, 1.305908236206044e+17, 1.305908236327922e+17, 1.305908236451364e+17, 1.305908236573242e+17, 1.305908236695119e+17, 1.305908236816998e+17, 1.305908236938876e+17, 1.305908237062317e+17, 1.305908237184195e+17, 1.305908237306074e+17, 1.305908237427951e+17, 1.305908237549829e+17, 1.305908237671708e+17, 1.305908237795148e+17, 1.305908237917027e+17, 1.305908238038904e+17, 1.305908238160783e+17, 1.305908238282661e+17, 1.305908238406102e+17, 1.305908238527981e+17, 1.305908238649857e+17, 1.305908238771736e+17, 1.305908238893614e+17, 1.305908239015493e+17, 1.305908239138934e+17, 1.305908239260812e+17, 1.305908239382691e+17, 1.305908239506131e+17, 1.305908239628009e+17, 1.305908239749887e+17, 1.305908239871766e+17, 1.305908239993644e+17, 1.305908240115521e+17, 1.305908240238963e+17, 1.30590824036084e+17, 1.305908240482719e+17, 1.305908240604596e+17, 1.305908240726476e+17, 1.305908240849916e+17, 1.305908240971794e+17, 1.305908241093673e+17, 1.305908241215551e+17, 1.305908241337428e+17, 1.305908241460869e+17, 1.305908241582748e+17, 1.305908241704626e+17, 1.305908241826504e+17, 1.305908241948383e+17, 1.30590824207026e+17, 1.305908242193701e+17, 1.305908242315579e+17, 1.305908242437458e+17, 1.305908242560897e+17, 1.305908242682778e+17, 1.305908242804655e+17, 1.305908242926533e+17, 1.305908243049974e+17, 1.305908243171852e+17, 1.305908243293731e+17, 1.305908243415608e+17, 1.305908243537486e+17, 1.305908243660927e+17, 1.305908243782806e+17, 1.305908243904685e+17, 1.305908244026563e+17, 1.30590824414844e+17, 1.305908244270318e+17, 1.305908244393759e+17, 1.305908244515636e+17, 1.305908244637516e+17, 1.305908244759395e+17, 1.305908244882834e+17, 1.305908245004713e+17, 1.305908245126591e+17, 1.30590824524847e+17, 1.305908245371909e+17, 1.305908245493788e+17, 1.305908245615666e+17, 1.305908245737545e+17, 1.305908245860986e+17, 1.305908245982863e+17, 1.305908246104742e+17, 1.305908246226619e+17, 1.305908246348498e+17, 1.305908246470376e+17, 1.305908246592253e+17, 1.305908246715695e+17, 1.305908246837573e+17, 1.305908246959452e+17, 1.30590824708133e+17, 1.305908247203208e+17, 1.305908247326648e+17, 1.305908247448526e+17, 1.305908247570406e+17, 1.305908247692283e+17, 1.305908247814162e+17, 1.30590824793604e+17, 1.305908248057917e+17, 1.305908248181358e+17, 1.305908248303236e+17, 1.305908248426678e+17, 1.305908248548556e+17, 1.305908248670435e+17, 1.305908248792312e+17, 1.30590824891419e+17, 1.305908249037631e+17, 1.30590824915951e+17, 1.305908249281388e+17, 1.305908249403265e+17, 1.305908249526706e+17, 1.305908249648585e+17, 1.305908249770463e+17, 1.30590824989234e+17, 1.305908250015782e+17, 1.30590825013766e+17, 1.305908250259538e+17, 1.305908250382979e+17, 1.305908250504858e+17, 1.305908250626735e+17, 1.305908250748613e+17, 1.305908250870492e+17, 1.30590825099237e+17, 1.305908251115811e+17, 1.305908251237688e+17, 1.305908251359566e+17, 1.305908251481446e+17, 1.305908251603324e+17, 1.305908251725202e+17, 1.305908251848643e+17, 1.30590825197052e+17, 1.305908252092399e+17, 1.305908252214277e+17, 1.305908252336156e+17, 1.305908252458034e+17, 1.305908252581475e+17, 1.305908252703352e+17, 1.30590825282523e+17, 1.305908252947109e+17, 1.305908253068987e+17, 1.305908253190865e+17, 1.305908253312744e+17, 1.305908253436184e+17, 1.305908253558062e+17, 1.30590825367994e+17, 1.305908253801819e+17, 1.305908253923697e+17, 1.305908254045574e+17, 1.305908254169016e+17, 1.305908254290894e+17, 1.305908254412773e+17, 1.305908254536212e+17, 1.305908254658092e+17, 1.305908254779969e+17, 1.30590825490341e+17, 1.305908255025288e+17, 1.305908255147167e+17, 1.305908255269044e+17, 1.305908255390922e+17, 1.305908255512801e+17, 1.305908255636242e+17, 1.305908255758121e+17, 1.305908255879999e+17, 1.305908256001876e+17, 1.305908256123756e+17, 1.305908256245633e+17, 1.305908256367511e+17, 1.305908256490952e+17, 1.305908256611267e+17, 1.305908256733146e+17, 1.305908256856586e+17, 1.305908256978464e+17, 1.305908257101905e+17, 1.305908257223785e+17, 1.305908257345661e+17, 1.30590825746754e+17, 1.305908257589418e+17, 1.305908257711296e+17, 1.305908257834738e+17, 1.305908257956614e+17, 1.305908258078495e+17, 1.305908258200372e+17, 1.305908258323813e+17, 1.305908258445691e+17, 1.305908258567569e+17, 1.305908258689448e+17, 1.305908258811324e+17, 1.305908258933203e+17, 1.305908259056644e+17, 1.305908259178523e+17, 1.305908259300401e+17, 1.305908259423841e+17, 1.30590825954572e+17, 1.305908259667598e+17, 1.305908259789476e+17, 1.305908259911355e+17, 1.305908260034796e+17, 1.305908260156673e+17, 1.305908260278551e+17, 1.30590826040043e+17, 1.305908260522308e+17, 1.305908260644186e+17, 1.305908260766063e+17, 1.305908260889505e+17, 1.305908261011383e+17, 1.305908261133261e+17, 1.30590826125514e+17, 1.305908261377018e+17, 1.305908261498897e+17, 1.305908261620774e+17, 1.305908261744215e+17, 1.305908261866094e+17, 1.305908261987972e+17, 1.305908262109851e+17, 1.305908262231727e+17, 1.305908262353605e+17, 1.305908262475484e+17, 1.305908262598925e+17, 1.305908262720804e+17, 1.305908262842682e+17, 1.305908262964559e+17, 1.305908263086437e+17, 1.305908263209879e+17, 1.305908263331757e+17, 1.305908263453635e+17, 1.305908263575514e+17, 1.305908263698953e+17, 1.305908263820833e+17, 1.305908263942711e+17, 1.305908264064589e+17, 1.305908264186467e+17, 1.305908264309907e+17, 1.305908264431785e+17, 1.305908264553663e+17, 1.305908264677105e+17, 1.305908264798982e+17, 1.305908264920861e+17, 1.305908265042739e+17, 1.30590826516618e+17, 1.305908265288058e+17, 1.305908265409935e+17, 1.305908265531814e+17, 1.305908265653693e+17, 1.305908265775571e+17, 1.305908265899012e+17, 1.30590826602089e+17, 1.305908266142767e+17, 1.305908266264645e+17, 1.305908266386524e+17, 1.305908266508402e+17, 1.305908266631844e+17, 1.305908266753722e+17, 1.305908266875599e+17, 1.305908266997478e+17, 1.305908267119356e+17, 1.305908267241235e+17, 1.305908267364675e+17, 1.305908267486554e+17, 1.305908267608433e+17, 1.305908267730309e+17, 1.305908267852188e+17, 1.305908267974066e+17, 1.305908268097507e+17, 1.305908268219384e+17, 1.305908268341263e+17, 1.305908268463142e+17, 1.30590826858502e+17, 1.305908268708461e+17, 1.305908268830339e+17, 1.305908268952218e+17, 1.305908269074095e+17, 1.305908269195973e+17, 1.305908269317852e+17, 1.30590826943973e+17, 1.305908269563171e+17, 1.305908269685048e+17, 1.305908269806927e+17, 1.305908269928805e+17, 1.305908270050683e+17, 1.305908270172562e+17, 1.30590827029444e+17, 1.30590827041788e+17, 1.305908270539758e+17, 1.305908270661637e+17, 1.305908270783515e+17, 1.305908270905393e+17, 1.305908271027272e+17, 1.305908271150711e+17, 1.305908271272591e+17, 1.305908271394469e+17, 1.305908271516347e+17, 1.305908271638226e+17, 1.305908271761665e+17, 1.305908271883544e+17, 1.305908272005421e+17, 1.3059082721273e+17, 1.305908272249179e+17, 1.305908272371057e+17, 1.305908272494497e+17, 1.305908272616375e+17, 1.305908272738254e+17, 1.305908272860132e+17, 1.305908272983572e+17, 1.305908273105452e+17, 1.305908273227329e+17, 1.305908273349208e+17, 1.305908273471086e+17, 1.305908273594527e+17, 1.305908273716404e+17, 1.305908273838284e+17, 1.305908273961723e+17, 1.305908274083602e+17, 1.305908274207043e+17, 1.305908274328922e+17, 1.305908274450799e+17, 1.305908274572677e+17, 1.305908274694556e+17, 1.305908274817996e+17, 1.305908274939875e+17, 1.305908275061752e+17, 1.30590827518363e+17, 1.305908275305509e+17, 1.30590827542895e+17, 1.305908275550828e+17, 1.305908275672705e+17, 1.305908275794584e+17, 1.305908275918025e+17, 1.305908276039904e+17, 1.305908276161782e+17, 1.305908276285222e+17, 1.3059082764071e+17, 1.305908276528978e+17, 1.305908276650857e+17, 1.305908276774298e+17, 1.305908276896177e+17, 1.305908277019616e+17, 1.305908277141495e+17, 1.305908277263373e+17, 1.305908277385252e+17, 1.30590827750713e+17, 1.305908277588381e+17, 1.305908277669633e+17, 1.305908277750886e+17, 1.305908277833701e+17, 1.305908277914953e+17, 1.305908277996205e+17, 1.305908278077457e+17, 1.305908278158708e+17, 1.30590827823996e+17, 1.305908278321212e+17, 1.305908278402465e+17, 1.30590827848528e+17, 1.305908278566532e+17, 1.305908278647784e+17, 1.305908278769663e+17, 1.30590827889154e+17, 1.305908279013418e+17, 1.305908279135297e+17, 1.305908279258738e+17, 1.305908279380616e+17, 1.305908279502493e+17, 1.305908279624372e+17, 1.305908279746252e+17, 1.305908279869692e+17, 1.30590827999157e+17, 1.305908280113448e+17, 1.305908280235327e+17, 1.305908280357204e+17, 1.305908280479082e+17, 1.305908280602523e+17, 1.305908280724402e+17, 1.305908280847843e+17, 1.30590828096972e+17, 1.305908281091598e+17, 1.305908281213476e+17, 1.305908281335355e+17, 1.305908281457234e+17, 1.305908281580675e+17, 1.305908281702552e+17, 1.30590828182443e+17, 1.305908281946309e+17, 1.305908282068187e+17, 1.305908282190065e+17, 1.305908282313505e+17, 1.305908282435384e+17, 1.305908282557262e+17, 1.30590828267914e+17, 1.305908282801019e+17, 1.305908282924458e+17, 1.305908283046337e+17, 1.305908283168215e+17, 1.305908283290094e+17, 1.305908283411972e+17, 1.305908283535412e+17, 1.305908283657292e+17, 1.305908283779169e+17, 1.305908283901048e+17, 1.305908284022926e+17, 1.305908284144803e+17, 1.305908284266683e+17, 1.305908284390122e+17, 1.305908284512001e+17, 1.305908284633879e+17, 1.305908284755757e+17, 1.305908284877636e+17, 1.305908285001076e+17, 1.305908285122954e+17, 1.305908285244832e+17, 1.305908285366711e+17, 1.305908285488589e+17, 1.305908285612031e+17, 1.305908285733908e+17, 1.305908285857349e+17, 1.305908285979227e+17, 1.305908286101105e+17, 1.305908286222984e+17, 1.305908286344861e+17, 1.30590828646674e+17, 1.305908286588618e+17, 1.305908286712059e+17, 1.305908286832374e+17, 1.305908286954253e+17, 1.305908287077693e+17, 1.305908287199571e+17, 1.305908287323013e+17, 1.305908287444891e+17, 1.305908287566769e+17, 1.305908287688646e+17, 1.305908287810524e+17, 1.305908287932403e+17, 1.305908288054282e+17, 1.30590828817616e+17, 1.305908288299601e+17, 1.305908288421478e+17, 1.305908288543357e+17, 1.305908288665235e+17, 1.305908288787113e+17, 1.305908288908992e+17, 1.30590828903087e+17, 1.30590828915431e+17, 1.305908289274627e+17, 1.305908289398067e+17, 1.305908289519945e+17, 1.305908289641823e+17, 1.305908289765265e+17, 1.305908289887142e+17, 1.305908290009021e+17, 1.305908290130899e+17, 1.305908290252777e+17, 1.305908290374655e+17, 1.305908290498097e+17, 1.305908290619974e+17, 1.305908290741852e+17, 1.305908290863731e+17, 1.305908290985609e+17, 1.305908291107487e+17, 1.305908291230927e+17, 1.305908291352805e+17, 1.305908291474684e+17, 1.305908291596562e+17, 1.305908291720004e+17, 1.305908291841882e+17, 1.305908291963759e+17, 1.305908292085638e+17, 1.305908292207515e+17, 1.305908292329394e+17, 1.305908292452835e+17, 1.305908292574714e+17, 1.305908292698153e+17, 1.305908292820032e+17, 1.30590829294191e+17, 1.305908293063789e+17, 1.305908293185667e+17, 1.305908293309107e+17, 1.305908293430986e+17, 1.305908293552864e+17, 1.305908293674743e+17, 1.305908293796621e+17, 1.305908293918497e+17, 1.305908294041939e+17, 1.305908294163817e+17, 1.305908294285695e+17, 1.305908294407574e+17, 1.305908294529452e+17, 1.305908294652892e+17, 1.305908294774771e+17, 1.305908294896649e+17, 1.305908295018527e+17, 1.305908295140406e+17, 1.305908295262284e+17, 1.305908295384161e+17, 1.305908295507603e+17, 1.305908295629481e+17, 1.305908295751359e+17, 1.305908295873236e+17, 1.305908295995116e+17, 1.305908296116993e+17, 1.305908296240435e+17, 1.305908296362313e+17, 1.305908296484191e+17, 1.30590829660607e+17, 1.305908296727946e+17, 1.305908296851388e+17, 1.305908296973266e+17, 1.305908297095144e+17, 1.305908297218586e+17, 1.305908297340463e+17, 1.305908297462342e+17, 1.30590829758422e+17, 1.305908297706098e+17, 1.305908297827976e+17, 1.305908297951418e+17, 1.305908298073295e+17, 1.305908298195173e+17, 1.305908298317052e+17, 1.305908298438929e+17, 1.305908298560808e+17, 1.305908298684248e+17, 1.305908298806127e+17, 1.305908298928005e+17, 1.305908299049883e+17, 1.305908299171762e+17, 1.305908299295203e+17, 1.30590829941708e+17},
			             {1.305907805993056e+17, 1.305907831082785e+17, 1.305907831164037e+17, 1.305907831245289e+17, 1.305907831326542e+17, 1.305907831489046e+17, 1.305907831570299e+17, 1.305907831651551e+17, 1.305907831734365e+17, 1.30590783189687e+17, 1.305907831978122e+17, 1.30590783890018e+17, 1.305907838979871e+17, 1.305907839143937e+17, 1.305907839225189e+17, 1.305907839306441e+17, 1.305907839387693e+17, 1.305907839468946e+17, 1.305907839550198e+17, 1.305907839714264e+17, 1.305907839795516e+17, 1.305907843540929e+17},
			             {1.305907806969646e+17, 1.305907846962894e+17},
			             {1.305907971789655e+17, 1.30590829941708e+17};
			mask_depths = {{0.5,  0.5, 10.4, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5, 10.4}, {0.5,  0.5, 10.4, 10.4}}, {{10.4,  10.4, 109.0, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 108.9}, {10.4, 108.9}, {10.4, 108.8}, {10.4, 108.7}, {10.4, 108.6}, {10.4, 108.5}, {10.4, 108.4}, {10.4, 108.4}, {10.4, 108.3}, {10.4, 108.3}, {10.4, 108.2}, {10.4, 108.2}, {10.4, 108.1}, {10.4, 108.1}, {10.4, 108.0}, {10.4, 107.9}, {10.4, 107.9}, {10.4, 107.8}, {10.4, 107.8}, {10.4, 107.7}, {10.4, 107.7}, {10.4, 107.6}, {10.4, 107.5}, {10.4, 107.5}, {10.4, 107.5}, {10.4, 107.4}, {10.4, 107.4}, {10.4, 107.4}, {10.4, 107.4}, {10.4, 107.3}, {10.4, 107.3}, {10.4, 107.3}, {10.4, 107.2}, {10.4, 107.2}, {10.4, 107.2}, {10.4, 107.2}, {10.4, 107.1}, {10.4, 107.1}, {10.4, 107.1}, {10.4, 107.1}, {10.4, 107.0}, {10.4, 107.0}, {10.4, 107.0}, {10.4, 107.0}, {10.4, 106.9}, {10.4, 106.9}, {10.4, 106.9}, {10.4, 106.9}, {10.4, 106.9}, {10.4, 106.8}, {10.4, 106.8}, {10.4, 106.8}, {10.4, 106.8}, {10.4, 106.8}, {10.4, 106.7}, {10.4, 106.7}, {10.4, 106.7}, {10.4, 106.7}, {10.4, 106.7}, {10.4, 106.6}, {10.4, 106.6}, {10.4, 106.6}, {10.4, 106.6}, {10.4, 106.6}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.5}, {10.4, 106.6}, {10.4, 106.6}, {10.4, 106.6}, {10.4, 106.7}, {10.4, 106.7}, {10.4, 106.8}, {10.4, 106.8}, {10.4, 106.8}, {10.4, 106.9}, {10.4, 106.9}, {10.4, 107.0}, {10.4, 107.0}, {10.4, 107.0}, {10.4, 107.1}, {10.4, 107.1}, {10.4, 107.2}, {10.4, 107.2}, {10.4, 107.2}, {10.4, 107.3}, {10.4, 107.3}, {10.4, 107.4}, {10.4, 107.4}, {10.4, 107.4}, {10.4, 107.5}, {10.4, 107.5}, {10.4, 107.6}, {10.4, 107.6}, {10.4, 107.7}, {10.4, 107.7}, {10.4, 107.7}, {10.4, 107.8}, {10.4, 107.8}, {10.4, 107.9}, {10.4, 107.9}, {10.4, 107.9}, {10.4, 108.0}, {10.4, 108.1}, {10.4, 108.1}, {10.4, 108.2}, {10.4, 108.3}, {10.4, 108.4}, {10.4, 108.5}, {10.4, 108.5}, {10.4, 108.5}, {10.4, 108.5}, {10.4, 108.5}, {10.4, 108.5}, {10.4, 108.6}, {10.4, 108.6}, {10.4, 108.7}, {10.4, 108.8}, {10.4, 108.9}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.1}, {10.4, 109.1}, {10.4, 109.1}, {10.4, 109.2}, {10.4, 109.2}, {10.4, 109.3}, {10.4, 109.3}, {10.4, 109.3}, {10.4, 109.4}, {10.4, 109.4}, {10.4, 110.0}, {10.4, 110.0}, {10.4, 110.0}, {10.4, 110.0}, {10.4, 110.0}, {10.4, 110.0}, {10.4, 110.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4,  10.4, 109.0, 109.0}}, {{10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4,  10.4, 109.0, 109.0}}, {{10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4,  10.4, 109.0, 109.0}}, {{10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4, 109.0}, {10.4,  10.4, 109.0, 109.0}}, {{41.6, 49.6}, {49.6}, {49.7}, {49.7}, {49.8}, {49.8}, {49.9}, {49.9}, {50.0}, {50.0}, {50.1}, {41.6}, {41.7}, {41.7}, {41.8}, {41.8}, {41.9}, {41.9}, {42.0}, {42.0}, {42.1}, {42.1, 50.1, 50.1}}, {{72.3, 80.3}, {72.3, 80.3}}, {{0.0, 9999.0}, {0.0, 9999.0}};
		}
	}
}
