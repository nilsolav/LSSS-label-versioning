netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 3;
			channels = 4;
			categories = 12;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  13.0, 13.0, 13.0;
			max_depth =  72.5, 71.8, 74.4;
			start_time = 129798778442470016, 129798778442470016, 129798771864344960;
			end_time = 129798778442470016, 129798778442470016, 129798778442470016;
			region_id = 1, 2, 3;
			region_name = "Layer1","Layer2","Layer3";
			region_provenance = "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "";
			region_category_names = "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12;
			region_type = analysis, analysis, analysis;
			channel_names = "18", "38", "200", "333";
			region_channels = 15, 15, 15;
			mask_times = {1.2979877844247e+17},
			             {1.2979877844247e+17},
			             {1.29798771864345e+17, 1.297987718763762e+17, 1.297987718884076e+17, 1.297987719004388e+17, 1.2979877191247e+17, 1.297987719245012e+17, 1.297987719365325e+17, 1.297987719485637e+17, 1.297987719607512e+17, 1.297987719727825e+17, 1.297987719848138e+17, 1.297987719968451e+17, 1.297987720088762e+17, 1.297987720209075e+17, 1.297987720329388e+17, 1.2979877204497e+17, 1.297987720570013e+17, 1.297987720690324e+17, 1.2979877208122e+17, 1.297987720932512e+17, 1.297987721052824e+17, 1.297987721173138e+17, 1.29798772129345e+17, 1.297987721413763e+17, 1.297987721534075e+17, 1.297987721654387e+17, 1.2979877217747e+17, 1.297987721896575e+17, 1.297987722016887e+17, 1.297987722137201e+17, 1.297987722257512e+17, 1.297987722377824e+17, 1.297987722498138e+17, 1.29798772261845e+17, 1.297987722738762e+17, 1.297987722860637e+17, 1.29798772298095e+17, 1.297987723101262e+17, 1.297987723221574e+17, 1.297987723341888e+17, 1.2979877234622e+17, 1.297987723582513e+17, 1.297987723702825e+17, 1.297987723823137e+17, 1.297987723943451e+17, 1.297987724065325e+17, 1.297987724185638e+17, 1.297987724305951e+17, 1.297987724426262e+17, 1.297987724546575e+17, 1.297987724666888e+17, 1.2979877247872e+17, 1.297987724907514e+17, 1.297987725027825e+17, 1.297987725148137e+17, 1.297987725270012e+17, 1.297987725390324e+17, 1.297987725510638e+17, 1.29798772563095e+17, 1.297987725751263e+17, 1.297987725871575e+17, 1.297987725991887e+17, 1.2979877261122e+17, 1.297987726232513e+17, 1.297987726354387e+17, 1.297987726474701e+17, 1.297987726595012e+17, 1.297987726715324e+17, 1.297987726835638e+17, 1.29798772695595e+17, 1.297987727076262e+17, 1.297987727196575e+17, 1.297987727316887e+17, 1.297987727437199e+17, 1.297987727559075e+17, 1.297987727679387e+17, 1.2979877277997e+17, 1.297987727920013e+17, 1.297987728040324e+17, 1.297987728160637e+17, 1.297987728280951e+17, 1.297987728401262e+17, 1.297987728523139e+17, 1.297987728643451e+17, 1.297987728763762e+17, 1.297987728884076e+17, 1.297987729004388e+17, 1.2979877291247e+17, 1.297987729245012e+17, 1.297987729365325e+17, 1.297987729485637e+17, 1.297987729605951e+17, 1.297987729727825e+17, 1.297987729848138e+17, 1.297987729968451e+17, 1.297987730088763e+17, 1.297987730209075e+17, 1.297987730329388e+17, 1.2979877304497e+17, 1.297987730570013e+17, 1.297987730690324e+17, 1.2979877308122e+17, 1.297987730932512e+17, 1.297987731052824e+17, 1.297987731173138e+17, 1.29798773129345e+17, 1.297987731413763e+17, 1.297987731534075e+17, 1.297987731654387e+17, 1.2979877317747e+17, 1.297987731896575e+17, 1.297987732016887e+17, 1.297987732137201e+17, 1.297987732257513e+17, 1.297987732377824e+17, 1.297987732498138e+17, 1.29798773261845e+17, 1.297987732738762e+17, 1.297987732859075e+17, 1.297987732979387e+17, 1.297987733101262e+17, 1.297987733221574e+17, 1.297987733341887e+17, 1.2979877334622e+17, 1.297987733582513e+17, 1.297987733702825e+17, 1.297987733823137e+17, 1.29798773394345e+17, 1.297987734063763e+17, 1.297987734185638e+17, 1.297987734305951e+17, 1.297987734426262e+17, 1.297987734546575e+17, 1.297987734666888e+17, 1.2979877347872e+17, 1.297987734907514e+17, 1.297987735027825e+17, 1.297987735148137e+17, 1.297987735268451e+17, 1.297987735390324e+17, 1.297987735510638e+17, 1.29798773563095e+17, 1.297987735751263e+17, 1.297987735871575e+17, 1.297987735991887e+17, 1.2979877361122e+17, 1.297987736232513e+17, 1.297987736352826e+17, 1.297987736474701e+17, 1.297987736595012e+17, 1.297987736715324e+17, 1.297987736835638e+17, 1.29798773695595e+17, 1.297987737076262e+17, 1.297987737196575e+17, 1.297987737316887e+17, 1.297987737437199e+17, 1.297987737559075e+17, 1.297987737679387e+17, 1.2979877377997e+17, 1.297987737920013e+17, 1.297987738040324e+17, 1.297987738160637e+17, 1.297987738280951e+17, 1.297987738401262e+17, 1.297987738521576e+17, 1.297987738641887e+17, 1.297987738763762e+17, 1.297987738884074e+17, 1.297987739004388e+17, 1.2979877391247e+17, 1.297987739245012e+17, 1.297987739365325e+17, 1.297987739485637e+17, 1.297987739605951e+17, 1.297987739727825e+17, 1.297987739848138e+17, 1.297987739968451e+17, 1.297987740088763e+17, 1.297987740209075e+17, 1.297987740329388e+17, 1.2979877404497e+17, 1.297987740570013e+17, 1.297987740690326e+17, 1.297987740810637e+17, 1.297987740932512e+17, 1.297987741052824e+17, 1.297987741173138e+17, 1.29798774129345e+17, 1.297987741413763e+17, 1.297987741534075e+17, 1.297987741654387e+17, 1.2979877417747e+17, 1.297987741895013e+17, 1.297987742015325e+17, 1.297987742137201e+17, 1.297987742257513e+17, 1.297987742377824e+17, 1.297987742498138e+17, 1.29798774261845e+17, 1.297987742738762e+17, 1.297987742859076e+17, 1.297987742979387e+17, 1.297987743101262e+17, 1.297987743221574e+17, 1.297987743341887e+17, 1.2979877434622e+17, 1.297987743582513e+17, 1.297987743702825e+17, 1.297987743823137e+17, 1.29798774394345e+17, 1.297987744063762e+17, 1.297987744184076e+17, 1.297987744305951e+17, 1.297987744426263e+17, 1.297987744546574e+17, 1.297987744666888e+17, 1.2979877447872e+17, 1.297987744907512e+17, 1.297987745027825e+17, 1.297987745148137e+17, 1.297987745268449e+17, 1.297987745390324e+17, 1.297987745510638e+17, 1.29798774563095e+17, 1.297987745751263e+17, 1.297987745871575e+17, 1.297987745991887e+17, 1.2979877461122e+17, 1.297987746232513e+17, 1.297987746352826e+17, 1.297987746473138e+17, 1.297987746595013e+17, 1.297987746715324e+17, 1.297987746835638e+17, 1.29798774695595e+17, 1.297987747076262e+17, 1.297987747196575e+17, 1.297987747316887e+17, 1.297987747437199e+17, 1.297987747557513e+17, 1.297987747679387e+17, 1.2979877477997e+17, 1.297987747920013e+17, 1.297987748040325e+17, 1.297987748160637e+17, 1.29798774828095e+17, 1.297987748401262e+17, 1.297987748521576e+17, 1.297987748641887e+17, 1.297987748763763e+17, 1.297987748884074e+17, 1.297987749004387e+17, 1.2979877491247e+17, 1.297987749245012e+17, 1.297987749365325e+17, 1.297987749485637e+17, 1.297987749605951e+17, 1.297987749726262e+17, 1.297987749848138e+17, 1.297987749968451e+17, 1.297987750088763e+17, 1.297987750209075e+17, 1.297987750329388e+17, 1.2979877504497e+17, 1.297987750570013e+17, 1.297987750690326e+17, 1.297987750810637e+17, 1.297987750932512e+17, 1.297987751052824e+17, 1.297987751173138e+17, 1.29798775129345e+17, 1.297987751413763e+17, 1.297987751534075e+17, 1.297987751654387e+17, 1.2979877517747e+17, 1.297987751895013e+17, 1.297987752015325e+17, 1.297987752137201e+17, 1.297987752257513e+17, 1.297987752377824e+17, 1.297987752498138e+17, 1.29798775261845e+17, 1.297987752738762e+17, 1.297987752859076e+17, 1.297987752979387e+17, 1.297987753099699e+17, 1.297987753221574e+17, 1.297987753341887e+17, 1.2979877534622e+17, 1.297987753582513e+17, 1.297987753702825e+17, 1.297987753823137e+17, 1.29798775394345e+17, 1.297987754063762e+17, 1.297987754184076e+17, 1.297987754304388e+17, 1.297987754426263e+17, 1.297987754546574e+17, 1.297987754666886e+17, 1.2979877547872e+17, 1.297987754907512e+17, 1.297987755027826e+17, 1.297987755148137e+17, 1.297987755268449e+17, 1.297987755388763e+17, 1.297987755510638e+17, 1.29798775563095e+17, 1.297987755751263e+17, 1.297987755871575e+17, 1.297987755991887e+17, 1.2979877561122e+17, 1.297987756232513e+17, 1.297987756352826e+17, 1.297987756473138e+17, 1.297987756595013e+17, 1.297987756715324e+17, 1.297987756835638e+17, 1.29798775695595e+17, 1.297987757076262e+17, 1.297987757196576e+17, 1.297987757316887e+17, 1.297987757437199e+17, 1.297987757557513e+17, 1.297987757677825e+17, 1.2979877577997e+17, 1.297987757920013e+17, 1.297987758040325e+17, 1.297987758160637e+17, 1.29798775828095e+17, 1.297987758401262e+17, 1.297987758521576e+17, 1.297987758641888e+17, 1.297987758763763e+17, 1.297987758884074e+17, 1.297987759004387e+17, 1.2979877591247e+17, 1.297987759245012e+17, 1.297987759365325e+17, 1.297987759485637e+17, 1.297987759605951e+17, 1.297987759726262e+17, 1.297987759846575e+17, 1.297987759968451e+17, 1.297987760088763e+17, 1.297987760209075e+17, 1.297987760329388e+17, 1.2979877604497e+17, 1.297987760570012e+17, 1.297987760690326e+17, 1.297987760810638e+17, 1.29798776093095e+17, 1.297987761052824e+17, 1.297987761173138e+17, 1.29798776129345e+17, 1.297987761413763e+17, 1.297987761534075e+17, 1.297987761654387e+17, 1.2979877617747e+17, 1.297987761895013e+17, 1.297987762015325e+17, 1.297987762135638e+17, 1.297987762257513e+17, 1.297987762377825e+17, 1.297987762498138e+17, 1.29798776261845e+17, 1.297987762738762e+17, 1.297987762859076e+17, 1.297987762979388e+17, 1.297987763099699e+17, 1.297987763220013e+17, 1.297987763341887e+17, 1.2979877634622e+17, 1.297987763582513e+17, 1.297987763702825e+17, 1.297987763823137e+17, 1.29798776394345e+17, 1.297987764063762e+17, 1.297987764184076e+17, 1.297987764304388e+17, 1.297987764426263e+17, 1.297987764546575e+17, 1.297987764666886e+17, 1.2979877647872e+17, 1.297987764907512e+17, 1.297987765027825e+17, 1.297987765148137e+17, 1.297987765268449e+17, 1.297987765388762e+17, 1.297987765509075e+17, 1.29798776563095e+17, 1.297987765751263e+17, 1.297987765871575e+17, 1.297987765991887e+17, 1.2979877661122e+17, 1.297987766232512e+17, 1.297987766352826e+17, 1.297987766473138e+17, 1.29798776659345e+17, 1.297987766715325e+17, 1.297987766835638e+17, 1.29798776695595e+17, 1.297987767076262e+17, 1.297987767196576e+17, 1.297987767316887e+17, 1.297987767437199e+17, 1.297987767557513e+17, 1.297987767677825e+17, 1.2979877677997e+17, 1.297987767920013e+17, 1.297987768040325e+17, 1.297987768160637e+17, 1.29798776828095e+17, 1.297987768401262e+17, 1.297987768521576e+17, 1.297987768641888e+17, 1.297987768762199e+17, 1.297987768882513e+17, 1.297987769004387e+17, 1.2979877691247e+17, 1.297987769245012e+17, 1.297987769365325e+17, 1.297987769485637e+17, 1.297987769605949e+17, 1.297987769726262e+17, 1.297987769846575e+17, 1.297987769966888e+17, 1.297987770088763e+17, 1.297987770209075e+17, 1.297987770329388e+17, 1.2979877704497e+17, 1.297987770570012e+17, 1.297987770690324e+17, 1.297987770810638e+17, 1.29798777093095e+17, 1.297987771051261e+17, 1.297987771173138e+17, 1.29798777129345e+17, 1.297987771413763e+17, 1.297987771534076e+17, 1.297987771654387e+17, 1.2979877717747e+17, 1.297987771895013e+17, 1.297987772015325e+17, 1.297987772135638e+17, 1.297987772257513e+17, 1.297987772377825e+17, 1.297987772498138e+17, 1.29798777261845e+17, 1.297987772738762e+17, 1.297987772859076e+17, 1.297987772979388e+17, 1.297987773099699e+17, 1.297987773220013e+17, 1.297987773340325e+17, 1.2979877734622e+17, 1.297987773582513e+17, 1.297987773702825e+17, 1.297987773823137e+17, 1.29798777394345e+17, 1.297987774063762e+17, 1.297987774184076e+17, 1.297987774304388e+17, 1.2979877744247e+17, 1.297987774545012e+17, 1.297987774666886e+17, 1.2979877747872e+17, 1.297987774907512e+17, 1.297987775027825e+17, 1.297987775148138e+17, 1.297987775268449e+17, 1.297987775388762e+17, 1.297987775509075e+17, 1.29798777563095e+17, 1.297987775751263e+17, 1.297987775871575e+17, 1.297987775991887e+17, 1.2979877761122e+17, 1.297987776232512e+17, 1.297987776352826e+17, 1.297987776473138e+17, 1.29798777659345e+17, 1.297987776715325e+17, 1.297987776835638e+17, 1.29798777695595e+17, 1.297987777076262e+17, 1.297987777196576e+17, 1.297987777316888e+17, 1.297987777437199e+17, 1.297987777557513e+17, 1.297987777677825e+17, 1.297987777798138e+17, 1.297987777920013e+17, 1.297987778040325e+17, 1.297987778160637e+17, 1.29798777828095e+17, 1.297987778401262e+17, 1.297987778521576e+17, 1.297987778641888e+17, 1.2979877787622e+17, 1.297987778882513e+17, 1.297987779004387e+17, 1.2979877791247e+17, 1.297987779245012e+17, 1.297987779365325e+17, 1.297987779485638e+17, 1.297987779605949e+17, 1.297987779726262e+17, 1.297987779846575e+17, 1.297987779966888e+17, 1.2979877800872e+17, 1.297987780209075e+17, 1.297987780329388e+17, 1.2979877804497e+17, 1.297987780570012e+17, 1.297987780690324e+17, 1.297987780810638e+17, 1.29798778093095e+17, 1.297987781051261e+17, 1.297987781173137e+17, 1.29798778129345e+17, 1.297987781413763e+17, 1.297987781534075e+17, 1.297987781654387e+17, 1.2979877817747e+17, 1.297987781895012e+17, 1.297987782015325e+17, 1.297987782135638e+17, 1.29798778225595e+17, 1.297987782377825e+17, 1.297987782498138e+17, 1.29798778261845e+17, 1.297987782738762e+17, 1.297987782859076e+17, 1.297987782979388e+17, 1.297987783099699e+17, 1.297987783220013e+17, 1.297987783340325e+17, 1.297987783460637e+17, 1.297987783582513e+17, 1.297987783702825e+17, 1.297987783823137e+17, 1.29798778394345e+17, 1.297987784063762e+17, 1.297987784184076e+17, 1.297987784304388e+17, 1.2979877844247e+17};
			mask_depths = {{}}, {{}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
