netcdf mask {
	:date_created = "20200810T140900";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200810T140900";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 22;
			channels = 6;
			categories = 132;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0, 21.2, 20.7, 19.9, 24.3, 19.2, 17.3, 18.8, 18.6, 27.2, 27.1, 35.5, 25.9, 28.9, 33.6, 28.8,  2.4, 63.1,  3.9, 64.3, 20.2, 38.6;
			max_depth =  75.0, 34.6, 34.5, 24.9, 31.2, 25.9, 31.7, 24.7, 34.7, 35.8, 34.7, 46.6, 38.8, 43.8, 37.8, 43.6,  2.8, 66.3,  4.1, 67.7, 22.5, 45.2;
			start_time = 131376810441888256, 131376817067200768, 131376811774388224, 131376811962669440, 131376812029857024, 131376812074388224, 131376812235169536, 131376812638607104, 131376812893294464, 131376818492669568, 131376819050169472, 131376825916732032, 131376827864700800, 131376828991419520, 131376829317981952, 131376829617200768, 131376828167981952, 131376827970794496, 131376832800794496, 131376825672513280, 131376821250638336, 131376832738294400;
			end_time = 131376832800794496, 131376817115638272, 131376811839544448, 131376811987044480, 131376812040169600, 131376812092825728, 131376812289232000, 131376812651419520, 131376812930325760, 131376818552669568, 131376819063607040, 131376825996107008, 131376827911888256, 131376829102044544, 131376829332513280, 131376829838138240, 131376828167981952, 131376828010638208, 131376832800794496, 131376825712982016, 131376821254857088, 131376832770638208;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22;
			region_name = "Layer1","Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "0", "0", "0", "0", "0", "0", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "6009", "6009", "6009", "6009", "6009", "6009", "5027", "5027", "5027", "5027", "5027", "5027", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "6009", "6009", "6009", "6009", "6009", "6009", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "6009", "6009", "6009", "6009", "6009", "6009", "1", "1", "1", "1", "1", "1", "6009", "6009", "6009", "6009", "6009", "6009", "0", "0", "0", "0", "0", "0", "1", "1", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63;
			mask_times = {1.313768104418883e+17, 1.313768104515758e+17, 1.313768104570446e+17, 1.313768104668883e+17, 1.313768104711071e+17, 1.31376810476732e+17, 1.313768104906382e+17, 1.31376810500482e+17, 1.313768105047007e+17, 1.313768105142321e+17, 1.313768105242319e+17, 1.313768105284507e+17, 1.31376810542982e+17, 1.313768105487633e+17, 1.31376810552982e+17, 1.313768105672008e+17, 1.313768105737633e+17, 1.313768105779821e+17, 1.313768105922007e+17, 1.313768105978257e+17, 1.313768106020444e+17, 1.313768106162633e+17, 1.31376810620482e+17, 1.313768106290757e+17, 1.313768106378257e+17, 1.313768106464195e+17, 1.31376810660482e+17, 1.313768106709508e+17, 1.313768106751695e+17, 1.313768106839195e+17, 1.313768106931382e+17, 1.313768107039195e+17, 1.313768107081382e+17, 1.313768107184507e+17, 1.31376810728607e+17, 1.313768107376695e+17, 1.313768107475133e+17, 1.31376810751732e+17, 1.313768107609508e+17, 1.313768107745445e+17, 1.313768107795444e+17, 1.31376810789232e+17, 1.313768107989194e+17, 1.313768108031382e+17, 1.313768108132945e+17, 1.313768108222008e+17, 1.31376810832357e+17, 1.313768108365757e+17, 1.313768108453257e+17, 1.313768108539195e+17, 1.313768108625133e+17, 1.313768108678258e+17, 1.313768108815757e+17, 1.313768108912632e+17, 1.31376810900482e+17, 1.31376810909857e+17, 1.31376810919857e+17, 1.313768109309508e+17, 1.313768109406383e+17, 1.313768109450132e+17, 1.313768109547008e+17, 1.31376810964857e+17, 1.313768109745445e+17, 1.313768109787633e+17, 1.313768109878257e+17, 1.313768109964195e+17, 1.31376811005482e+17, 1.313768110153258e+17, 1.313768110251695e+17, 1.313768110301695e+17, 1.313768110407945e+17, 1.313768110506383e+17, 1.313768110548571e+17, 1.31376811063607e+17, 1.313768110740756e+17, 1.313768110839195e+17, 1.313768110895444e+17, 1.31376811099232e+17, 1.31376811103607e+17, 1.313768111142319e+17, 1.313768111239195e+17, 1.313768111281382e+17, 1.313768111373571e+17, 1.313768111459508e+17, 1.313768111559507e+17, 1.313768111656383e+17, 1.31376811169857e+17, 1.31376811179232e+17, 1.313768111878258e+17, 1.313768111965757e+17, 1.313768112059507e+17, 1.31376811215482e+17, 1.313768112253257e+17, 1.313768112314195e+17, 1.313768112412632e+17, 1.313768112457944e+17, 1.313768112543882e+17, 1.31376811262982e+17, 1.313768112725133e+17, 1.31376811282982e+17, 1.313768112926694e+17, 1.31376811302982e+17, 1.313768113072008e+17, 1.313768113159507e+17, 1.313768113245445e+17, 1.31376811333607e+17, 1.31376811342982e+17, 1.31376811352982e+17, 1.313768113626694e+17, 1.313768113718883e+17, 1.313768113762633e+17, 1.313768113851694e+17, 1.313768113939195e+17, 1.313768114045445e+17, 1.313768114150132e+17, 1.313768114247008e+17, 1.313768114295444e+17, 1.313768114395444e+17, 1.313768114493883e+17, 1.31376811453607e+17, 1.31376811459232e+17, 1.313768114725133e+17, 1.313768114831383e+17, 1.313768114873571e+17, 1.313768115022007e+17, 1.313768115068883e+17, 1.313768115164195e+17, 1.313768115264196e+17, 1.313768115362632e+17, 1.31376811546107e+17, 1.313768115559507e+17, 1.313768115614195e+17, 1.313768115714195e+17, 1.313768115811071e+17, 1.313768115915757e+17, 1.313768115957944e+17, 1.313768116051695e+17, 1.313768116153257e+17, 1.313768116251695e+17, 1.313768116293882e+17, 1.313768116382944e+17, 1.313768116475132e+17, 1.313768116573569e+17, 1.313768116675132e+17, 1.313768116776695e+17, 1.31376811682357e+17, 1.313768116914195e+17, 1.313768117015757e+17, 1.313768117114195e+17, 1.313768117173569e+17, 1.313768117272008e+17, 1.31376811732357e+17, 1.31376811742982e+17, 1.313768117528257e+17, 1.313768117570445e+17, 1.313768117657944e+17, 1.313768117743882e+17, 1.31376811788607e+17, 1.313768117951694e+17, 1.31376811804857e+17, 1.31376811810482e+17, 1.313768118206382e+17, 1.313768118256383e+17, 1.313768118395444e+17, 1.31376811844857e+17, 1.313768118547008e+17, 1.31376811863607e+17, 1.313768118728257e+17, 1.313768118772008e+17, 1.313768118857944e+17, 1.313768118943884e+17, 1.31376811902982e+17, 1.31376811911732e+17, 1.31376811920482e+17, 1.313768119297009e+17, 1.313768119339195e+17, 1.313768119395444e+17, 1.313768119487633e+17, 1.313768119626694e+17, 1.31376811972357e+17, 1.313768119770445e+17, 1.313768119870445e+17, 1.313768119912632e+17, 1.31376812005482e+17, 1.313768120114195e+17, 1.313768120156383e+17, 1.31376812029857e+17, 1.313768120359508e+17, 1.313768120401696e+17, 1.313768120500133e+17, 1.313768120606382e+17, 1.313768120701695e+17, 1.313768120743882e+17, 1.31376812088607e+17, 1.313768120928257e+17, 1.313768121018883e+17, 1.313768121114195e+17, 1.313768121200132e+17, 1.31376812128607e+17, 1.313768121381382e+17, 1.313768121470445e+17, 1.313768121556383e+17, 1.313768121645444e+17, 1.313768121736069e+17, 1.313768121823571e+17, 1.313768121926696e+17, 1.313768122025133e+17, 1.313768122131382e+17, 1.313768122190757e+17, 1.313768122287633e+17, 1.313768122351695e+17, 1.31376812244857e+17, 1.313768122490757e+17, 1.313768122576695e+17, 1.313768122636069e+17, 1.313768122734508e+17, 1.313768122790757e+17, 1.31376812289232e+17, 1.31376812293607e+17, 1.313768123037632e+17, 1.313768123131383e+17, 1.313768123228257e+17, 1.313768123332945e+17, 1.313768123382944e+17, 1.31376812348607e+17, 1.313768123584507e+17, 1.313768123681382e+17, 1.31376812372357e+17, 1.313768123809508e+17, 1.313768123950134e+17, 1.31376812399857e+17, 1.313768124097007e+17, 1.313768124187633e+17, 1.31376812428607e+17, 1.313768124384507e+17, 1.313768124426694e+17, 1.313768124567319e+17, 1.313768124625133e+17, 1.313768124711071e+17, 1.313768124797007e+17, 1.313768124884507e+17, 1.313768124970446e+17, 1.313768125106382e+17, 1.313768125150132e+17, 1.313768125289194e+17, 1.313768125334508e+17, 1.313768125443882e+17, 1.313768125534508e+17, 1.313768125625133e+17, 1.313768125717321e+17, 1.313768125814195e+17, 1.313768125912634e+17, 1.313768125962633e+17, 1.31376812606107e+17, 1.313768126104819e+17, 1.31376812619857e+17, 1.313768126284508e+17, 1.313768126386071e+17, 1.313768126428257e+17, 1.313768126514195e+17, 1.313768126609508e+17, 1.313768126701696e+17, 1.313768126806382e+17, 1.313768126903258e+17, 1.313768126957944e+17, 1.313768127059507e+17, 1.31376812716107e+17, 1.313768127207945e+17, 1.313768127309508e+17, 1.313768127407945e+17, 1.313768127453257e+17, 1.313768127539195e+17, 1.313768127626696e+17, 1.313768127712632e+17, 1.313768127811069e+17, 1.313768127907945e+17, 1.313768127964195e+17, 1.313768128062633e+17, 1.31376812810482e+17, 1.31376812815482e+17, 1.313768128284507e+17, 1.313768128370445e+17, 1.313768128457946e+17, 1.313768128557944e+17, 1.313768128656381e+17, 1.31376812869857e+17, 1.31376812878607e+17, 1.31376812883607e+17, 1.313768128932945e+17, 1.313768129075132e+17, 1.31376812916107e+17, 1.313768129247008e+17, 1.313768129303258e+17, 1.313768129442321e+17, 1.31376812950482e+17, 1.313768129609507e+17, 1.313768129651695e+17, 1.313768129740758e+17, 1.313768129828257e+17, 1.313768129914195e+17, 1.313768130056383e+17, 1.31376813015482e+17, 1.313768130197007e+17, 1.31376813030482e+17, 1.313768130407945e+17, 1.313768130500133e+17, 1.313768130557944e+17, 1.313768130656383e+17, 1.31376813069857e+17, 1.31376813078607e+17, 1.313768130872008e+17, 1.313768130975132e+17, 1.31376813101732e+17, 1.313768131190757e+17, 1.313768131234508e+17, 1.313768131325133e+17, 1.313768131411071e+17, 1.313768131553257e+17, 1.313768131648571e+17, 1.313768131747007e+17, 1.313768131843882e+17, 1.31376813188607e+17, 1.313768131973569e+17, 1.313768132114195e+17, 1.313768132157946e+17, 1.313768132293883e+17, 1.313768132342321e+17, 1.31376813242982e+17, 1.313768132525133e+17, 1.313768132620445e+17, 1.313768132712632e+17, 1.313768132853257e+17, 1.313768132906383e+17, 1.313768133006382e+17, 1.31376813304857e+17, 1.313768133193883e+17, 1.313768133236069e+17, 1.313768133334508e+17, 1.313768133431382e+17, 1.31376813352982e+17, 1.313768133578258e+17, 1.313768133675132e+17, 1.313768133773571e+17, 1.313768133815758e+17, 1.31376813400482e+17, 1.313768134064195e+17, 1.313768134162633e+17, 1.313768134211071e+17, 1.313768134297007e+17, 1.313768134437632e+17, 1.313768134489196e+17, 1.313768134575133e+17, 1.313768134662633e+17, 1.31376813479857e+17, 1.313768134884508e+17, 1.313768134972008e+17, 1.313768135062633e+17, 1.31376813516107e+17, 1.313768135206383e+17, 1.31376813533607e+17, 1.313768135378258e+17, 1.313768135468883e+17, 1.31376813556732e+17, 1.313768135665757e+17, 1.313768135709508e+17, 1.313768135806382e+17, 1.313768135907945e+17, 1.313768136003258e+17, 1.313768136100133e+17, 1.313768136142321e+17, 1.31376813622982e+17, 1.313768136370445e+17, 1.313768136412632e+17, 1.313768136520445e+17, 1.313768136617321e+17, 1.31376813666732e+17, 1.31376813676732e+17, 1.313768136864195e+17, 1.313768136914195e+17, 1.313768137012632e+17, 1.313768137109508e+17, 1.313768137151695e+17, 1.313768137245444e+17, 1.313768137342319e+17, 1.313768137384508e+17, 1.313768137526694e+17, 1.313768137568882e+17, 1.31376813769857e+17, 1.313768137800133e+17, 1.313768137897007e+17, 1.313768137989196e+17, 1.313768138032945e+17, 1.313768138125133e+17, 1.313768138211069e+17, 1.31376813829857e+17, 1.313768138437632e+17, 1.31376813847982e+17, 1.31376813856732e+17, 1.313768138707945e+17, 1.313768138765757e+17, 1.313768138865757e+17, 1.313768138951695e+17, 1.313768139037632e+17, 1.313768139145445e+17, 1.313768139187633e+17, 1.31376813929232e+17, 1.313768139334508e+17, 1.313768139390757e+17, 1.313768139539196e+17, 1.313768139626694e+17, 1.31376813971732e+17, 1.313768139806383e+17, 1.313768139906382e+17, 1.313768140004819e+17, 1.313768140056383e+17, 1.31376814014857e+17, 1.313768140245445e+17, 1.313768140297007e+17, 1.313768140382945e+17, 1.313768140468883e+17, 1.313768140522008e+17, 1.31376814065482e+17, 1.313768140742321e+17, 1.313768140828257e+17, 1.313768140972008e+17, 1.31376814101732e+17, 1.313768141109507e+17, 1.313768141207945e+17, 1.313768141250132e+17, 1.313768141342321e+17, 1.313768141442319e+17, 1.313768141545445e+17, 1.31376814160482e+17, 1.313768141648571e+17, 1.313768141734508e+17, 1.313768141875132e+17, 1.31376814193607e+17, 1.313768141978257e+17, 1.313768142065757e+17, 1.31376814216107e+17, 1.31376814226107e+17, 1.313768142357946e+17, 1.313768142459507e+17, 1.313768142518883e+17, 1.31376814256107e+17, 1.31376814266107e+17, 1.313768142765757e+17, 1.313768142864195e+17, 1.313768142965757e+17, 1.313768143056383e+17, 1.31376814309857e+17, 1.313768143245445e+17, 1.31376814329857e+17, 1.313768143395446e+17, 1.313768143447008e+17, 1.313768143543882e+17, 1.313768143642319e+17, 1.313768143690757e+17, 1.313768143789194e+17, 1.31376814388607e+17, 1.313768143928257e+17, 1.313768144022008e+17, 1.313768144126696e+17, 1.313768144168883e+17, 1.313768144256383e+17, 1.313768144311069e+17, 1.31376814444857e+17, 1.313768144542319e+17, 1.313768144584507e+17, 1.313768144672008e+17, 1.313768144757944e+17, 1.313768144843882e+17, 1.313768144934508e+17, 1.31376814502982e+17, 1.313768145126694e+17, 1.313768145168882e+17, 1.313768145256383e+17, 1.313768145303258e+17, 1.313768145431383e+17, 1.313768145518883e+17, 1.31376814566732e+17, 1.313768145715757e+17, 1.313768145822008e+17, 1.313768145864195e+17, 1.313768145920444e+17, 1.31376814604857e+17, 1.313768146145444e+17, 1.313768146242319e+17, 1.313768146284508e+17, 1.313768146370445e+17, 1.313768146457946e+17, 1.313768146547007e+17, 1.31376814664857e+17, 1.313768146745445e+17, 1.313768146790757e+17, 1.313768146889196e+17, 1.31376814698607e+17, 1.313768147037632e+17, 1.313768147132945e+17, 1.31376814722982e+17, 1.313768147272008e+17, 1.313768147365757e+17, 1.313768147473571e+17, 1.313768147526696e+17, 1.313768147625133e+17, 1.31376814772357e+17, 1.313768147773571e+17, 1.313768147872008e+17, 1.313768147970446e+17, 1.313768148018883e+17, 1.31376814810482e+17, 1.313768148201696e+17, 1.313768148309507e+17, 1.313768148351694e+17, 1.313768148406382e+17, 1.313768148545445e+17, 1.313768148642319e+17, 1.313768148739195e+17, 1.31376814878607e+17, 1.313768148872008e+17, 1.313768149007945e+17, 1.313768149064196e+17, 1.313768149106383e+17, 1.313768149253257e+17, 1.313768149301696e+17, 1.313768149403258e+17, 1.313768149500132e+17, 1.313768149557944e+17, 1.313768149659508e+17, 1.313768149701696e+17, 1.313768149789196e+17, 1.313768149882944e+17, 1.313768149982945e+17, 1.313768150081382e+17, 1.31376815012357e+17, 1.313768150225133e+17, 1.313768150325132e+17, 1.31376815036732e+17, 1.313768150462633e+17, 1.31376815055482e+17, 1.313768150656383e+17, 1.31376815069857e+17, 1.313768150839195e+17, 1.313768150893883e+17, 1.313768150995446e+17, 1.313768151093883e+17, 1.31376815119232e+17, 1.313768151234508e+17, 1.313768151322007e+17, 1.313768151415758e+17, 1.313768151514195e+17, 1.31376815161732e+17, 1.313768151672008e+17, 1.313768151714195e+17, 1.313768151865757e+17, 1.313768151907945e+17, 1.313768151995444e+17, 1.313768152087633e+17, 1.313768152184507e+17, 1.313768152231383e+17, 1.31376815231732e+17, 1.313768152412632e+17, 1.313768152511071e+17, 1.313768152553257e+17, 1.313768152640756e+17, 1.313768152726696e+17, 1.313768152812632e+17, 1.31376815290482e+17, 1.313768153001696e+17, 1.313768153103258e+17, 1.313768153147008e+17, 1.313768153281382e+17, 1.31376815332357e+17, 1.313768153411069e+17, 1.313768153551694e+17, 1.313768153607945e+17, 1.313768153701695e+17, 1.313768153745445e+17, 1.313768153875132e+17, 1.313768153918883e+17, 1.313768154014195e+17, 1.313768154109508e+17, 1.313768154207945e+17, 1.31376815426732e+17, 1.313768154309508e+17, 1.313768154395444e+17, 1.313768154539195e+17, 1.313768154597007e+17, 1.313768154695446e+17, 1.313768154743882e+17, 1.313768154845445e+17, 1.313768154942319e+17, 1.313768154989196e+17, 1.313768155095444e+17, 1.313768155137632e+17, 1.313768155228257e+17, 1.313768155320445e+17, 1.313768155412632e+17, 1.313768155511071e+17, 1.313768155553257e+17, 1.313768155645445e+17, 1.313768155743882e+17, 1.31376815578607e+17, 1.313768155873571e+17, 1.31376815596107e+17, 1.313768156053257e+17, 1.313768156148571e+17, 1.313768156251695e+17, 1.313768156293883e+17, 1.313768156381382e+17, 1.313768156515757e+17, 1.31376815656107e+17, 1.313768156651695e+17, 1.313768156750132e+17, 1.313768156797007e+17, 1.313768156882945e+17, 1.313768156984507e+17, 1.313768157081382e+17, 1.31376815712357e+17, 1.313768157214195e+17, 1.313768157312632e+17, 1.31376815735482e+17, 1.313768157495444e+17, 1.313768157545445e+17, 1.313768157642321e+17, 1.313768157684508e+17, 1.313768157742319e+17, 1.313768157840756e+17, 1.313768157981382e+17, 1.31376815802357e+17, 1.313768158111071e+17, 1.313768158211069e+17, 1.313768158309508e+17, 1.313768158353258e+17, 1.313768158447007e+17, 1.313768158537632e+17, 1.313768158632945e+17, 1.313768158675133e+17, 1.313768158765757e+17, 1.313768158862633e+17, 1.313768158959507e+17, 1.313768159001695e+17, 1.313768159107945e+17, 1.31376815919857e+17, 1.313768159290757e+17, 1.31376815939232e+17, 1.313768159495444e+17, 1.313768159550132e+17, 1.31376815959232e+17, 1.31376815969857e+17, 1.313768159795444e+17, 1.313768159862632e+17, 1.31376815996107e+17, 1.313768160018883e+17, 1.313768160112632e+17, 1.313768160211069e+17, 1.313768160268882e+17, 1.313768160311071e+17, 1.313768160412634e+17, 1.313768160511069e+17, 1.313768160559508e+17, 1.313768160700133e+17, 1.313768160756383e+17, 1.31376816079857e+17, 1.313768160939195e+17, 1.31376816098607e+17, 1.313768161078257e+17, 1.313768161168882e+17, 1.313768161214195e+17, 1.313768161311071e+17, 1.313768161409508e+17, 1.313768161506383e+17, 1.313768161564195e+17, 1.31376816166107e+17, 1.313768161703258e+17, 1.313768161801695e+17, 1.313768161900133e+17, 1.313768161951695e+17, 1.313768162043882e+17, 1.313768162142319e+17, 1.313768162190757e+17, 1.313768162289196e+17, 1.31376816238607e+17, 1.313768162443882e+17, 1.313768162545445e+17, 1.313768162587633e+17, 1.313768162678258e+17, 1.313768162776695e+17, 1.313768162875132e+17, 1.31376816291732e+17, 1.313768163003258e+17, 1.31376816309232e+17, 1.31376816319232e+17, 1.313768163297007e+17, 1.313768163357946e+17, 1.31376816345482e+17, 1.31376816349857e+17, 1.313768163584508e+17, 1.31376816367982e+17, 1.313768163781382e+17, 1.313768163882945e+17, 1.313768163981382e+17, 1.31376816402982e+17, 1.313768164134508e+17, 1.313768164232945e+17, 1.31376816432982e+17, 1.313768164389196e+17, 1.31376816448607e+17, 1.313768164547008e+17, 1.313768164651695e+17, 1.313768164693882e+17, 1.31376816479232e+17, 1.313768164890757e+17, 1.313768164989196e+17, 1.313768165045444e+17, 1.313768165140758e+17, 1.313768165239195e+17, 1.313768165281382e+17, 1.313768165372008e+17, 1.313768165475132e+17, 1.313768165573571e+17, 1.31376816562357e+17, 1.313768165720444e+17, 1.313768165811069e+17, 1.313768165872008e+17, 1.313768165968882e+17, 1.313768166011069e+17, 1.313768166097007e+17, 1.31376816620482e+17, 1.313768166301695e+17, 1.31376816636107e+17, 1.313768166451695e+17, 1.313768166543882e+17, 1.31376816658607e+17, 1.313768166676695e+17, 1.313768166776695e+17, 1.313768166820444e+17, 1.313768166904819e+17, 1.31376816699232e+17, 1.313768167097007e+17, 1.313768167143882e+17, 1.313768167237632e+17, 1.313768167334508e+17, 1.313768167437632e+17, 1.313768167482945e+17, 1.313768167576695e+17, 1.313768167662632e+17, 1.313768167750132e+17, 1.313768167850132e+17, 1.31376816789232e+17, 1.313768167981382e+17, 1.313768168078258e+17, 1.313768168176695e+17, 1.313768168232945e+17, 1.313768168318883e+17, 1.313768168412632e+17, 1.313768168518883e+17, 1.31376816856107e+17, 1.31376816865482e+17, 1.313768168747008e+17, 1.313768168836069e+17, 1.313768168922007e+17, 1.31376816901732e+17, 1.313768169131383e+17, 1.31376816922982e+17, 1.313768169328257e+17, 1.313768169425133e+17, 1.313768169475132e+17, 1.313768169564195e+17, 1.313768169664196e+17, 1.313768169706382e+17, 1.313768169795444e+17, 1.313768169889196e+17, 1.313768169989196e+17, 1.313768170087633e+17, 1.313768170140758e+17, 1.313768170240758e+17, 1.313768170284508e+17, 1.313768170381382e+17, 1.313768170484508e+17, 1.313768170528257e+17, 1.31376817062982e+17, 1.313768170672008e+17, 1.313768170768882e+17, 1.313768170873571e+17, 1.313768170928257e+17, 1.313768171026696e+17, 1.313768171068883e+17, 1.313768171156383e+17, 1.313768171289194e+17, 1.313768171331383e+17, 1.313768171440758e+17, 1.313768171537632e+17, 1.313768171584508e+17, 1.313768171670445e+17, 1.313768171772008e+17, 1.313768171868882e+17, 1.313768171911069e+17, 1.313768172000132e+17, 1.313768172090757e+17, 1.313768172195444e+17, 1.313768172237632e+17, 1.31376817229232e+17, 1.313768172420444e+17, 1.313768172511069e+17, 1.313768172601695e+17, 1.313768172703258e+17, 1.313768172809508e+17, 1.313768172851694e+17, 1.313768172993883e+17, 1.313768173053257e+17, 1.313768173153258e+17, 1.313768173207945e+17, 1.313768173312632e+17, 1.31376817335482e+17, 1.313768173412632e+17, 1.313768173557946e+17, 1.313768173612632e+17, 1.313768173711071e+17, 1.313768173753258e+17, 1.313768173893883e+17, 1.313768173950132e+17, 1.313768174051695e+17, 1.313768174103256e+17, 1.313768174200132e+17, 1.313768174242321e+17, 1.31376817432982e+17, 1.31376817442357e+17, 1.313768174518883e+17, 1.313768174611071e+17, 1.313768174697007e+17, 1.313768174790757e+17, 1.313768174887631e+17, 1.313768174984507e+17, 1.313768175034508e+17, 1.313768175125133e+17, 1.313768175222007e+17, 1.313768175275132e+17, 1.313768175376695e+17, 1.313768175475132e+17, 1.313768175532946e+17, 1.313768175637632e+17, 1.313768175679821e+17, 1.313768175809508e+17, 1.313768175900133e+17, 1.313768176000133e+17, 1.31376817609857e+17, 1.313768176150132e+17, 1.31376817624857e+17, 1.313768176347008e+17, 1.313768176404819e+17, 1.313768176509508e+17, 1.313768176557944e+17, 1.313768176656383e+17, 1.31376817669857e+17, 1.31376817678607e+17, 1.313768176887633e+17, 1.313768176931383e+17, 1.31376817702982e+17, 1.313768177132945e+17, 1.313768177175133e+17, 1.313768177262632e+17, 1.31376817734857e+17, 1.313768177434508e+17, 1.313768177575133e+17, 1.313768177632945e+17, 1.313768177675132e+17, 1.313768177809507e+17, 1.313768177851695e+17, 1.313768177945445e+17, 1.313768178045444e+17, 1.313768178147008e+17, 1.313768178204819e+17, 1.31376817830482e+17, 1.313768178347008e+17, 1.313768178434508e+17, 1.313768178532945e+17, 1.313768178626696e+17, 1.31376817871732e+17, 1.313768178759508e+17, 1.313768178847007e+17, 1.313768178940758e+17, 1.313768178982945e+17, 1.313768179118883e+17, 1.313768179178258e+17, 1.313768179268883e+17, 1.313768179311069e+17, 1.313768179407945e+17, 1.313768179504819e+17, 1.313768179601695e+17, 1.31376817966107e+17, 1.313768179757944e+17, 1.313768179800132e+17, 1.313768179887633e+17, 1.313768179984507e+17, 1.31376818002982e+17, 1.313768180134508e+17, 1.313768180232945e+17, 1.313768180284508e+17, 1.313768180381382e+17, 1.313768180487633e+17, 1.313768180587633e+17, 1.313768180634508e+17, 1.313768180720445e+17, 1.31376818081732e+17, 1.313768180914195e+17, 1.313768180956381e+17, 1.313768181042319e+17, 1.313768181184508e+17, 1.313768181231383e+17, 1.313768181322007e+17, 1.313768181407945e+17, 1.313768181500133e+17, 1.313768181600132e+17, 1.31376818170482e+17, 1.313768181803258e+17, 1.313768181859507e+17, 1.313768181951695e+17, 1.313768181995444e+17, 1.313768182082945e+17, 1.313768182168882e+17, 1.313768182256383e+17, 1.313768182347008e+17, 1.313768182443882e+17, 1.313768182542319e+17, 1.313768182584507e+17, 1.313768182682945e+17, 1.31376818277982e+17, 1.313768182876695e+17, 1.313768182918883e+17, 1.313768183006383e+17, 1.313768183101695e+17, 1.313768183200133e+17, 1.313768183295444e+17, 1.31376818339232e+17, 1.313768183434508e+17, 1.313768183528257e+17, 1.313768183626696e+17, 1.313768183668883e+17, 1.313768183765757e+17, 1.313768183865757e+17, 1.313768183907945e+17, 1.313768183995446e+17, 1.313768184087633e+17, 1.31376818419232e+17, 1.313768184290757e+17, 1.313768184332945e+17, 1.313768184389194e+17, 1.31376818453607e+17, 1.313768184632945e+17, 1.31376818467982e+17, 1.313768184778257e+17, 1.313768184875132e+17, 1.313768184926696e+17, 1.313768185026694e+17, 1.313768185068882e+17, 1.31376818515482e+17, 1.31376818524857e+17, 1.31376818534857e+17, 1.313768185390757e+17, 1.313768185526696e+17, 1.313768185575133e+17, 1.313768185670445e+17, 1.313768185714195e+17, 1.313768185854821e+17, 1.313768185901695e+17, 1.313768186001696e+17, 1.313768186100132e+17, 1.31376818614857e+17, 1.313768186245445e+17, 1.313768186343882e+17, 1.313768186401696e+17, 1.313768186500133e+17, 1.313768186547008e+17, 1.313768186651695e+17, 1.31376818674857e+17, 1.313768186793882e+17, 1.31376818689857e+17, 1.313768186940756e+17, 1.313768187037632e+17, 1.313768187140756e+17, 1.313768187195444e+17, 1.313768187237632e+17, 1.313768187378257e+17, 1.313768187432945e+17, 1.313768187536069e+17, 1.313768187590757e+17, 1.313768187682945e+17, 1.313768187725133e+17, 1.31376818786732e+17, 1.313768187920445e+17, 1.313768188014195e+17, 1.313768188112632e+17, 1.313768188156383e+17, 1.313768188328257e+17, 1.313768188372008e+17, 1.313768188457944e+17, 1.313768188600133e+17, 1.313768188659507e+17, 1.313768188757946e+17, 1.313768188800132e+17, 1.31376818889232e+17, 1.313768188978258e+17, 1.313768189064196e+17, 1.313768189165757e+17, 1.313768189259507e+17, 1.313768189301695e+17, 1.313768189395444e+17, 1.313768189489196e+17, 1.313768189587633e+17, 1.31376818968607e+17, 1.313768189743882e+17, 1.313768189840758e+17, 1.313768189887633e+17, 1.313768190025133e+17, 1.31376819006732e+17, 1.31376819016732e+17, 1.313768190265757e+17, 1.313768190307945e+17, 1.313768190409507e+17, 1.313768190501695e+17, 1.313768190593883e+17, 1.31376819063607e+17, 1.313768190728257e+17, 1.313768190814195e+17, 1.313768190900132e+17, 1.313768190995444e+17, 1.313768191097007e+17, 1.313768191200133e+17, 1.31376819129232e+17, 1.313768191334508e+17, 1.313768191422007e+17, 1.313768191507945e+17, 1.313768191607945e+17, 1.313768191709508e+17, 1.313768191751694e+17, 1.313768191842319e+17, 1.313768191928257e+17, 1.313768192025133e+17, 1.313768192073569e+17, 1.313768192159507e+17, 1.31376819225482e+17, 1.313768192353257e+17, 1.313768192395444e+17, 1.313768192482945e+17, 1.313768192570445e+17, 1.313768192678258e+17, 1.313768192776695e+17, 1.313768192831383e+17, 1.313768192873571e+17, 1.313768193015757e+17, 1.313768193057944e+17, 1.31376819314857e+17, 1.313768193253257e+17, 1.313768193297007e+17, 1.313768193384508e+17, 1.313768193489194e+17, 1.313768193587633e+17, 1.31376819363607e+17, 1.313768193737632e+17, 1.31376819378607e+17, 1.313768193882944e+17, 1.31376819397982e+17, 1.313768194039195e+17, 1.31376819413607e+17, 1.313768194178258e+17, 1.313768194322007e+17, 1.31376819436732e+17, 1.313768194470445e+17, 1.313768194512634e+17, 1.313768194600132e+17, 1.313768194690757e+17, 1.313768194781382e+17, 1.313768194884508e+17, 1.313768194928257e+17, 1.313768195032945e+17, 1.313768195075132e+17, 1.313768195215758e+17, 1.313768195264195e+17, 1.313768195370445e+17, 1.313768195412632e+17, 1.313768195500132e+17, 1.313768195673571e+17, 1.31376819572982e+17, 1.313768195826696e+17, 1.313768195925132e+17, 1.313768195973569e+17, 1.313768196068883e+17, 1.313768196165757e+17, 1.313768196211069e+17, 1.313768196311071e+17, 1.313768196409508e+17, 1.313768196475133e+17, 1.31376819651732e+17, 1.31376819660482e+17, 1.31376819669232e+17, 1.313768196789196e+17, 1.313768196887633e+17, 1.31376819692982e+17, 1.313768197026696e+17, 1.313768197125133e+17, 1.31376819716732e+17, 1.31376819725482e+17, 1.313768197356383e+17, 1.313768197459507e+17, 1.313768197507945e+17, 1.313768197609508e+17, 1.313768197651695e+17, 1.313768197739195e+17, 1.313768197825133e+17, 1.313768197920445e+17, 1.313768198020444e+17, 1.313768198111069e+17, 1.313768198159507e+17, 1.313768198253258e+17, 1.313768198351695e+17, 1.313768198393883e+17, 1.313768198481382e+17, 1.313768198590757e+17, 1.313768198647007e+17, 1.313768198745445e+17, 1.313768198809508e+17, 1.313768198901695e+17, 1.313768198943882e+17, 1.313768199036069e+17, 1.313768199128257e+17, 1.313768199225133e+17, 1.31376819926732e+17, 1.313768199362633e+17, 1.313768199462633e+17, 1.313768199553257e+17, 1.313768199597007e+17, 1.313768199689196e+17, 1.313768199784508e+17, 1.313768199881382e+17, 1.31376819992357e+17, 1.313768200015758e+17, 1.31376820011732e+17, 1.313768200209508e+17, 1.313768200253258e+17, 1.313768200350134e+17, 1.313768200450132e+17, 1.313768200497007e+17, 1.313768200582945e+17, 1.313768200682945e+17, 1.313768200725132e+17, 1.313768200870445e+17, 1.313768200920445e+17, 1.313768201020445e+17, 1.313768201062633e+17, 1.313768201150132e+17, 1.313768201243882e+17, 1.313768201297007e+17, 1.313768201431383e+17, 1.313768201482945e+17, 1.313768201582945e+17, 1.313768201681382e+17, 1.313768201725133e+17, 1.313768201820445e+17, 1.313768201917321e+17, 1.31376820196107e+17, 1.313768202047008e+17, 1.313768202132945e+17, 1.313768202220445e+17, 1.313768202325133e+17, 1.313768202422008e+17, 1.313768202464196e+17, 1.313768202562633e+17, 1.313768202659507e+17, 1.313768202701696e+17, 1.313768202787633e+17, 1.313768202875132e+17, 1.313768202973571e+17, 1.313768203072008e+17, 1.313768203125133e+17, 1.313768203167319e+17, 1.313768203222007e+17, 1.313768203318883e+17, 1.313768203411071e+17, 1.313768203507945e+17, 1.313768203550132e+17, 1.313768203637633e+17, 1.313768203731382e+17, 1.31376820382982e+17, 1.313768203926694e+17, 1.313768203975132e+17, 1.313768204072008e+17, 1.313768204170445e+17, 1.31376820421732e+17, 1.31376820431732e+17, 1.313768204414195e+17, 1.31376820446732e+17, 1.313768204565757e+17, 1.313768204607945e+17, 1.31376820469857e+17, 1.31376820479857e+17, 1.313768204897007e+17, 1.313768204950132e+17, 1.313768205051695e+17, 1.313768205150132e+17, 1.313768205242319e+17, 1.313768205334508e+17, 1.313768205376695e+17, 1.313768205518883e+17, 1.313768205575132e+17, 1.313768205617321e+17, 1.313768205704819e+17, 1.313768205797007e+17, 1.313768205887633e+17, 1.31376820598607e+17, 1.313768206034508e+17, 1.313768206125133e+17, 1.31376820622357e+17, 1.313768206272008e+17, 1.313768206372008e+17, 1.313768206462633e+17, 1.31376820650482e+17, 1.31376820659232e+17, 1.313768206651695e+17, 1.313768206787631e+17, 1.313768206873571e+17, 1.313768206972008e+17, 1.313768207014195e+17, 1.31376820710482e+17, 1.313768207207945e+17, 1.313768207306383e+17, 1.313768207368882e+17, 1.313768207411071e+17, 1.313768207553257e+17, 1.313768207614195e+17, 1.313768207656381e+17, 1.31376820782982e+17, 1.313768207873571e+17, 1.313768207975133e+17, 1.313768208073569e+17, 1.31376820811732e+17, 1.313768208214195e+17, 1.313768208257944e+17, 1.313768208314195e+17, 1.313768208454821e+17, 1.313768208501695e+17, 1.313768208631383e+17, 1.313768208676695e+17, 1.313768208768882e+17, 1.313768208862633e+17, 1.31376820899232e+17, 1.313768209086071e+17, 1.313768209187633e+17, 1.313768209284507e+17, 1.313768209332945e+17, 1.31376820942982e+17, 1.313768209472008e+17, 1.313768209601695e+17, 1.31376820966107e+17, 1.313768209759507e+17, 1.313768209803258e+17, 1.313768209895444e+17, 1.313768209995444e+17, 1.313768210037632e+17, 1.313768210125133e+17, 1.31376821021732e+17, 1.31376821026107e+17, 1.313768210401695e+17, 1.313768210493882e+17, 1.313768210545445e+17, 1.313768210645444e+17, 1.31376821069232e+17, 1.313768210790757e+17, 1.313768210887633e+17, 1.313768210932945e+17, 1.31376821102982e+17, 1.313768211128257e+17, 1.313768211187633e+17, 1.313768211290758e+17, 1.313768211332945e+17, 1.313768211387633e+17, 1.313768211484507e+17, 1.313768211570445e+17, 1.313768211656383e+17, 1.313768211743882e+17, 1.313768211836069e+17, 1.313768211937632e+17, 1.313768211979821e+17, 1.313768212072008e+17, 1.313768212165757e+17, 1.313768212265757e+17, 1.313768212362633e+17, 1.313768212414195e+17, 1.313768212506383e+17, 1.313768212548571e+17, 1.313768212684508e+17, 1.313768212743882e+17, 1.313768212840758e+17, 1.313768212893883e+17, 1.31376821298607e+17, 1.313768213082945e+17, 1.313768213128257e+17, 1.313768213222007e+17, 1.313768213320445e+17, 1.313768213417321e+17, 1.313768213479821e+17, 1.313768213578257e+17, 1.313768213631383e+17, 1.313768213726696e+17, 1.313768213768883e+17, 1.31376821390482e+17, 1.31376821396732e+17, 1.313768214065757e+17, 1.313768214125133e+17, 1.31376821416732e+17, 1.313768214303258e+17, 1.31376821439857e+17, 1.31376821446107e+17, 1.313768214503258e+17, 1.313768214600132e+17, 1.313768214687633e+17, 1.313768214773571e+17, 1.313768214864195e+17, 1.313768214950132e+17, 1.313768215090757e+17, 1.313768215132945e+17, 1.313768215220444e+17, 1.313768215311069e+17, 1.31376821541732e+17, 1.313768215459508e+17, 1.313768215589196e+17, 1.313768215650132e+17, 1.31376821574857e+17, 1.313768215797007e+17, 1.313768215897007e+17, 1.313768215995444e+17, 1.313768216051695e+17, 1.313768216143882e+17, 1.31376821618607e+17, 1.313768216276695e+17, 1.313768216362633e+17, 1.313768216462633e+17, 1.31376821650482e+17, 1.313768216595444e+17, 1.313768216693883e+17, 1.31376821673607e+17, 1.31376821682357e+17, 1.313768216926694e+17, 1.313768216968882e+17, 1.313768217031383e+17, 1.313768217175132e+17, 1.313768217231382e+17, 1.31376821732982e+17, 1.313768217372008e+17, 1.313768217457946e+17, 1.313768217545445e+17, 1.313768217650132e+17, 1.313768217707945e+17, 1.313768217750132e+17, 1.313768217897007e+17, 1.313768217950132e+17, 1.31376821799232e+17, 1.31376821807982e+17, 1.313768218175132e+17, 1.313768218265757e+17, 1.313768218351695e+17, 1.313768218439195e+17, 1.31376821854857e+17, 1.313768218647008e+17, 1.313768218745445e+17, 1.313768218801695e+17, 1.313768218900133e+17, 1.313768218942319e+17, 1.313768218998569e+17, 1.313768219126694e+17, 1.313768219214195e+17, 1.313768219303258e+17, 1.313768219397007e+17, 1.313768219495444e+17, 1.313768219543882e+17, 1.31376821962982e+17, 1.313768219720444e+17, 1.313768219814195e+17, 1.313768219870445e+17, 1.313768219968882e+17, 1.313768220011071e+17, 1.31376822009857e+17, 1.313768220184508e+17, 1.313768220281382e+17, 1.313768220378258e+17, 1.31376822042357e+17, 1.313768220520445e+17, 1.313768220562633e+17, 1.313768220650132e+17, 1.313768220739195e+17, 1.313768220839195e+17, 1.313768220881382e+17, 1.31376822102982e+17, 1.313768221089196e+17, 1.313768221131382e+17, 1.313768221218883e+17, 1.313768221314195e+17, 1.31376822141732e+17, 1.313768221459507e+17, 1.31376822155482e+17, 1.313768221642321e+17, 1.313768221742321e+17, 1.313768221784507e+17, 1.313768221875132e+17, 1.313768221976695e+17, 1.313768222018883e+17, 1.31376822210482e+17, 1.313768222250132e+17, 1.31376822229232e+17, 1.313768222379821e+17, 1.313768222470445e+17, 1.313768222568882e+17, 1.313768222665757e+17, 1.313768222725133e+17, 1.313768222825133e+17, 1.31376822292357e+17, 1.313768223025133e+17, 1.313768223073571e+17, 1.313768223162633e+17, 1.313768223262632e+17, 1.31376822330482e+17, 1.31376822339232e+17, 1.313768223490757e+17, 1.313768223532945e+17, 1.313768223620444e+17, 1.313768223711071e+17, 1.313768223812634e+17, 1.313768223909508e+17, 1.313768223951695e+17, 1.313768224059507e+17, 1.313768224107945e+17, 1.313768224203258e+17, 1.313768224301695e+17, 1.313768224403258e+17, 1.313768224495444e+17, 1.313768224543882e+17, 1.313768224650132e+17, 1.313768224747008e+17, 1.313768224795446e+17, 1.313768224895444e+17, 1.313768224937632e+17, 1.313768225028257e+17, 1.313768225126696e+17, 1.31376822522357e+17, 1.313768225276695e+17, 1.313768225370445e+17, 1.313768225468882e+17, 1.31376822551732e+17, 1.313768225603258e+17, 1.313768225689196e+17, 1.313768225779821e+17, 1.313768225865757e+17, 1.313768225951695e+17, 1.313768226093882e+17, 1.31376822619232e+17, 1.31376822628607e+17, 1.313768226382945e+17, 1.313768226426694e+17, 1.313768226520445e+17, 1.313768226620445e+17, 1.313768226726694e+17, 1.313768226781382e+17, 1.31376822682357e+17, 1.313768226911071e+17, 1.313768227006382e+17, 1.313768227097007e+17, 1.313768227197007e+17, 1.313768227239195e+17, 1.313768227337633e+17, 1.313768227443882e+17, 1.31376822748607e+17, 1.313768227543882e+17, 1.313768227672008e+17, 1.313768227759507e+17, 1.313768227898569e+17, 1.313768227990757e+17, 1.313768228087633e+17, 1.31376822812982e+17, 1.313768228220444e+17, 1.313768228315757e+17, 1.313768228368883e+17, 1.31376822846732e+17, 1.313768228509508e+17, 1.313768228651695e+17, 1.313768228711069e+17, 1.31376822875482e+17, 1.313768228889194e+17, 1.313768228943882e+17, 1.313768229040756e+17, 1.313768229082944e+17, 1.313768229176695e+17, 1.313768229279821e+17, 1.31376822932357e+17, 1.313768229426694e+17, 1.313768229525133e+17, 1.31376822958607e+17, 1.313768229676695e+17, 1.313768229768882e+17, 1.313768229865757e+17, 1.313768229907945e+17, 1.31376823000482e+17, 1.313768230101695e+17, 1.313768230143882e+17, 1.31376823022982e+17, 1.31376823031732e+17, 1.313768230407945e+17, 1.313768230504819e+17, 1.313768230562633e+17, 1.31376823060482e+17, 1.313768230656381e+17, 1.31376823079857e+17, 1.313768230840758e+17, 1.313768230934508e+17, 1.313768231032945e+17, 1.31376823108607e+17, 1.313768231182945e+17, 1.313768231245445e+17, 1.313768231342319e+17, 1.313768231387633e+17, 1.31376823148607e+17, 1.313768231582945e+17, 1.313768231631383e+17, 1.313768231732945e+17, 1.313768231831383e+17, 1.313768231897007e+17, 1.313768231939195e+17, 1.313768232028257e+17, 1.313768232114195e+17, 1.313768232201695e+17, 1.313768232297007e+17, 1.313768232406382e+17, 1.31376823244857e+17, 1.313768232593883e+17, 1.313768232657944e+17, 1.313768232701695e+17, 1.313768232797009e+17, 1.313768232887633e+17, 1.313768232973571e+17, 1.313768233059507e+17, 1.313768233145445e+17, 1.313768233195444e+17, 1.313768233325133e+17, 1.313768233412632e+17, 1.313768233507945e+17, 1.313768233606382e+17, 1.313768233709508e+17, 1.31376823376107e+17, 1.313768233857944e+17, 1.313768233956383e+17, 1.313768234001695e+17, 1.313768234109508e+17, 1.313768234204819e+17, 1.313768234262633e+17, 1.31376823430482e+17, 1.313768234445445e+17, 1.313768234506382e+17, 1.31376823454857e+17, 1.313768234609508e+17, 1.313768234745445e+17, 1.313768234843884e+17, 1.31376823488607e+17, 1.313768234981382e+17, 1.313768235070445e+17, 1.31376823516107e+17, 1.313768235247008e+17, 1.313768235345445e+17, 1.313768235443882e+17, 1.313768235542321e+17, 1.31376823559232e+17, 1.313768235693883e+17, 1.31376823579857e+17, 1.313768235840758e+17, 1.313768235931383e+17, 1.313768236031382e+17, 1.313768236128257e+17, 1.31376823617982e+17, 1.31376823626732e+17, 1.313768236353257e+17, 1.313768236459507e+17, 1.313768236501695e+17, 1.313768236593883e+17, 1.313768236690757e+17, 1.313768236787633e+17, 1.31376823682982e+17, 1.31376823691732e+17, 1.313768237028257e+17, 1.313768237072008e+17, 1.313768237157946e+17, 1.313768237245445e+17, 1.313768237347008e+17, 1.313768237397007e+17, 1.313768237493883e+17, 1.313768237539195e+17, 1.31376823763607e+17, 1.313768237734508e+17, 1.313768237782944e+17, 1.31376823787982e+17, 1.313768237976695e+17, 1.313768238025133e+17, 1.31376823812357e+17, 1.313768238222008e+17, 1.313768238270445e+17, 1.313768238370445e+17, 1.31376823846732e+17, 1.313768238514195e+17, 1.313768238612632e+17, 1.31376823865482e+17, 1.313768238756383e+17, 1.313768238848571e+17, 1.313768238893883e+17, 1.313768238990757e+17, 1.313768239089194e+17, 1.313768239139195e+17, 1.313768239245445e+17, 1.313768239287633e+17, 1.313768239382945e+17, 1.313768239484507e+17, 1.313768239575132e+17, 1.313768239628257e+17, 1.313768239717321e+17, 1.313768239807945e+17, 1.313768239906382e+17, 1.313768239948571e+17, 1.313768240042319e+17, 1.31376824013607e+17, 1.313768240232945e+17, 1.313768240331383e+17, 1.313768240373571e+17, 1.31376824046732e+17, 1.313768240556383e+17, 1.31376824065482e+17, 1.313768240697007e+17, 1.31376824079232e+17, 1.31376824088607e+17, 1.313768240984507e+17, 1.313768241039195e+17, 1.313768241136069e+17, 1.313768241178257e+17, 1.313768241265757e+17, 1.313768241409508e+17, 1.313768241451694e+17, 1.313768241542319e+17, 1.313768241643882e+17, 1.313768241689194e+17, 1.313768241775132e+17, 1.313768241922008e+17, 1.313768241965757e+17, 1.313768242100132e+17, 1.313768242142321e+17, 1.313768242243884e+17, 1.313768242342321e+17, 1.313768242395446e+17, 1.313768242489194e+17, 1.313768242587633e+17, 1.31376824264857e+17, 1.313768242745445e+17, 1.313768242787633e+17, 1.313768242887633e+17, 1.31376824298607e+17, 1.31376824308607e+17, 1.313768243147007e+17, 1.313768243189194e+17, 1.31376824327982e+17, 1.313768243365757e+17, 1.313768243468882e+17, 1.31376824356732e+17, 1.313768243622008e+17, 1.313768243718883e+17, 1.313768243815757e+17, 1.313768243872008e+17, 1.313768243968883e+17, 1.313768244011071e+17, 1.313768244097007e+17, 1.313768244248571e+17, 1.313768244301695e+17, 1.31376824439857e+17, 1.313768244440756e+17, 1.313768244528257e+17, 1.31376824462357e+17, 1.313768244722008e+17, 1.313768244764196e+17, 1.313768244937632e+17, 1.313768244982945e+17, 1.313768245082944e+17, 1.313768245181382e+17, 1.31376824522982e+17, 1.313768245326694e+17, 1.31376824542357e+17, 1.313768245465757e+17, 1.313768245551694e+17, 1.313768245653257e+17, 1.313768245695446e+17, 1.31376824579232e+17, 1.313768245893883e+17, 1.313768245956383e+17, 1.313768246053257e+17, 1.313768246095446e+17, 1.313768246181382e+17, 1.313768246315758e+17, 1.313768246359507e+17, 1.313768246453258e+17, 1.313768246550132e+17, 1.31376824659232e+17, 1.313768246678258e+17, 1.313768246765757e+17, 1.313768246857944e+17, 1.313768246957946e+17, 1.313768247056383e+17, 1.313768247106382e+17, 1.313768247197007e+17, 1.313768247295444e+17, 1.313768247340758e+17, 1.313768247432945e+17, 1.313768247531382e+17, 1.313768247578258e+17, 1.313768247670445e+17, 1.313768247770445e+17, 1.313768247862633e+17, 1.313768247970445e+17, 1.313768248031382e+17, 1.31376824812982e+17, 1.31376824817982e+17, 1.31376824827982e+17, 1.313768248322007e+17, 1.313768248415758e+17, 1.313768248512632e+17, 1.313768248559507e+17, 1.313768248647008e+17, 1.31376824874857e+17, 1.313768248839195e+17, 1.313768248882945e+17, 1.313768248968883e+17, 1.313768249018883e+17, 1.313768249167319e+17, 1.313768249265757e+17, 1.313768249309508e+17, 1.313768249395444e+17, 1.313768249481382e+17, 1.313768249543882e+17, 1.313768249689196e+17, 1.313768249731382e+17, 1.313768249873571e+17, 1.313768249925133e+17, 1.313768250020445e+17, 1.313768250072008e+17, 1.313768250114195e+17, 1.313768250200132e+17, 1.313768250250132e+17, 1.31376825039232e+17, 1.313768250489196e+17, 1.313768250556383e+17, 1.31376825059857e+17, 1.31376825068607e+17, 1.313768250772008e+17, 1.313768250857946e+17, 1.313768250957944e+17, 1.31376825106107e+17, 1.313768251103258e+17, 1.313768251190757e+17, 1.313768251276695e+17, 1.313768251362633e+17, 1.31376825151732e+17, 1.313768251562633e+17, 1.313768251651695e+17, 1.313768251750132e+17, 1.31376825179232e+17, 1.313768251881382e+17, 1.31376825196732e+17, 1.313768252053257e+17, 1.313768252109508e+17, 1.313768252243884e+17, 1.313768252339195e+17, 1.313768252381382e+17, 1.31376825246732e+17, 1.313768252559508e+17, 1.313768252651695e+17, 1.313768252750132e+17, 1.31376825279232e+17, 1.31376825288607e+17, 1.31376825298607e+17, 1.313768253082945e+17, 1.313768253139195e+17, 1.313768253231382e+17, 1.313768253325133e+17, 1.313768253373571e+17, 1.31376825346732e+17, 1.313768253553257e+17, 1.31376825364857e+17, 1.313768253750132e+17, 1.313768253856383e+17, 1.313768253901696e+17, 1.313768253990757e+17, 1.313768254089196e+17, 1.313768254131383e+17, 1.313768254218883e+17, 1.31376825430482e+17, 1.313768254409508e+17, 1.313768254451694e+17, 1.31376825455482e+17, 1.313768254653257e+17, 1.313768254697007e+17, 1.313768254790757e+17, 1.313768254889196e+17, 1.313768254931382e+17, 1.313768255018883e+17, 1.313768255112632e+17, 1.31376825520482e+17, 1.313768255301695e+17, 1.313768255343882e+17, 1.313768255431382e+17, 1.313768255534508e+17, 1.313768255632946e+17, 1.313768255682945e+17, 1.313768255784508e+17, 1.31376825587982e+17, 1.313768255968882e+17, 1.313768256070445e+17, 1.31376825612357e+17, 1.313768256214195e+17, 1.313768256311069e+17, 1.313768256353257e+17, 1.313768256440758e+17, 1.313768256531383e+17, 1.313768256620444e+17, 1.313768256725133e+17, 1.313768256778257e+17, 1.313768256875132e+17, 1.313768256975133e+17, 1.31376825703607e+17, 1.31376825712982e+17, 1.313768257172008e+17, 1.313768257265757e+17, 1.313768257359508e+17, 1.313768257457944e+17, 1.313768257500133e+17, 1.313768257587633e+17, 1.313768257679821e+17, 1.313768257765757e+17, 1.313768257862633e+17, 1.313768257962633e+17, 1.313768258004819e+17, 1.313768258097007e+17, 1.313768258189194e+17, 1.313768258289196e+17, 1.313768258331383e+17, 1.31376825841732e+17, 1.31376825851732e+17, 1.313768258559507e+17, 1.313768258645445e+17, 1.313768258753257e+17, 1.313768258795444e+17, 1.313768258882945e+17, 1.313768258939195e+17, 1.313768259081382e+17, 1.31376825916732e+17, 1.313768259253258e+17, 1.313768259343882e+17, 1.31376825942982e+17, 1.313768259518883e+17, 1.313768259615757e+17, 1.313768259657944e+17, 1.313768259801696e+17, 1.313768259857944e+17, 1.31376825996107e+17, 1.313768260014195e+17, 1.313768260111071e+17, 1.313768260153257e+17, 1.313768260239195e+17, 1.313768260331383e+17, 1.31376826042982e+17, 1.313768260522007e+17, 1.313768260568882e+17, 1.313768260665757e+17, 1.313768260762633e+17, 1.31376826080482e+17, 1.313768260893883e+17, 1.313768260990758e+17, 1.313768261032945e+17, 1.313768261173571e+17, 1.313768261231382e+17, 1.313768261334508e+17, 1.313768261382944e+17, 1.313768261484508e+17, 1.313768261526696e+17, 1.313768261612632e+17, 1.313768261715757e+17, 1.313768261759507e+17, 1.313768261889196e+17, 1.313768261943882e+17, 1.313768262042321e+17, 1.313768262112632e+17, 1.31376826215482e+17, 1.313768262240756e+17, 1.313768262331382e+17, 1.31376826242982e+17, 1.313768262528257e+17, 1.313768262578258e+17, 1.313768262675132e+17, 1.313768262772008e+17, 1.313768262820445e+17, 1.313768262925133e+17, 1.31376826296732e+17, 1.313768263057944e+17, 1.313768263156383e+17, 1.313768263215757e+17, 1.313768263320445e+17, 1.313768263376695e+17, 1.313768263475132e+17, 1.31376826351732e+17, 1.313768263612632e+17, 1.313768263712632e+17, 1.31376826375482e+17, 1.313768263842319e+17, 1.313768263943882e+17, 1.313768264040758e+17, 1.313768264139195e+17, 1.313768264187633e+17, 1.313768264284508e+17, 1.313768264382945e+17, 1.313768264437633e+17, 1.313768264534508e+17, 1.313768264576695e+17, 1.313768264706382e+17, 1.313768264751695e+17, 1.313768264853257e+17, 1.313768264895444e+17, 1.313768264981382e+17, 1.313768265122008e+17, 1.31376826518607e+17, 1.313768265282945e+17, 1.313768265325133e+17, 1.31376826541732e+17, 1.313768265515757e+17, 1.313768265620445e+17, 1.313768265711071e+17, 1.313768265753258e+17, 1.313768265901695e+17, 1.313768265954821e+17, 1.313768265997007e+17, 1.313768266082945e+17, 1.313768266170445e+17, 1.313768266265757e+17, 1.31376826636107e+17, 1.313768266464196e+17, 1.31376826656732e+17, 1.313768266664195e+17, 1.313768266706382e+17, 1.31376826679232e+17, 1.31376826692982e+17, 1.313768267026696e+17, 1.313768267081382e+17, 1.313768267173569e+17, 1.313768267264195e+17, 1.313768267306382e+17, 1.313768267393883e+17, 1.313768267490757e+17, 1.313768267589196e+17, 1.313768267686071e+17, 1.313768267737632e+17, 1.313768267829819e+17, 1.313768267928257e+17, 1.313768267976695e+17, 1.313768268070445e+17, 1.31376826819232e+17, 1.313768268282945e+17, 1.313768268382944e+17, 1.313768268426696e+17, 1.313768268512632e+17, 1.313768268653257e+17, 1.313768268706383e+17, 1.31376826880482e+17, 1.31376826885482e+17, 1.313768268953257e+17, 1.313768269043882e+17, 1.31376826909232e+17, 1.313768269187633e+17, 1.313768269284508e+17, 1.313768269328257e+17, 1.313768269418883e+17, 1.313768269512632e+17, 1.313768269611071e+17, 1.313768269657944e+17, 1.313768269751695e+17, 1.313768269850132e+17, 1.313768269953258e+17, 1.313768269995444e+17, 1.313768270082945e+17, 1.313768270168882e+17, 1.31376827025482e+17, 1.313768270395444e+17, 1.313768270437633e+17, 1.313768270528257e+17, 1.313768270620445e+17, 1.313768270712632e+17, 1.31376827075482e+17, 1.313768270900133e+17, 1.313768270956383e+17, 1.31376827099857e+17, 1.31376827108607e+17, 1.313768271172008e+17, 1.313768271276695e+17, 1.313768271373571e+17, 1.31376827143607e+17, 1.313768271536069e+17, 1.313768271579821e+17, 1.313768271689196e+17, 1.313768271790757e+17, 1.313768271834508e+17, 1.31376827192982e+17, 1.313768272026694e+17, 1.313768272068883e+17, 1.31376827216107e+17, 1.31376827226107e+17, 1.313768272357946e+17, 1.31376827241732e+17, 1.313768272507945e+17, 1.313768272606383e+17, 1.31376827266732e+17, 1.313768272765757e+17, 1.313768272814195e+17, 1.313768272906382e+17, 1.313768273003258e+17, 1.313768273095444e+17, 1.313768273137632e+17, 1.31376827323607e+17, 1.313768273332945e+17, 1.313768273437632e+17, 1.31376827347982e+17, 1.313768273570445e+17, 1.313768273673569e+17, 1.313768273773571e+17, 1.313768273872008e+17, 1.313768273968883e+17, 1.31376827406732e+17, 1.313768274115757e+17, 1.313768274217321e+17, 1.313768274265757e+17, 1.313768274356383e+17, 1.31376827449857e+17, 1.313768274542319e+17, 1.313768274637632e+17, 1.31376827473607e+17, 1.313768274778257e+17, 1.313768274834508e+17, 1.313768274976695e+17, 1.313768275072008e+17, 1.313768275114195e+17, 1.313768275207945e+17, 1.313768275309508e+17, 1.313768275351695e+17, 1.313768275437633e+17, 1.313768275532945e+17, 1.31376827562357e+17, 1.313768275723571e+17, 1.313768275765757e+17, 1.313768275822007e+17, 1.313768275950132e+17, 1.313768276036069e+17, 1.31376827612357e+17, 1.313768276209508e+17, 1.313768276306383e+17, 1.31376827640482e+17, 1.313768276447008e+17, 1.31376827659232e+17, 1.313768276643882e+17, 1.313768276734508e+17, 1.313768276776695e+17, 1.313768276864195e+17, 1.313768276956383e+17, 1.313768277048571e+17, 1.313768277090757e+17, 1.313768277262633e+17, 1.313768277318883e+17, 1.31376827741732e+17, 1.313768277473571e+17, 1.313768277576695e+17, 1.313768277618883e+17, 1.31376827772357e+17, 1.313768277765757e+17, 1.313768277901695e+17, 1.313768277943882e+17, 1.313768278087633e+17, 1.313768278137632e+17, 1.313768278225133e+17, 1.313768278328257e+17, 1.313768278370445e+17, 1.313768278457946e+17, 1.313768278550132e+17, 1.313768278647008e+17, 1.313768278743882e+17, 1.313768278787633e+17, 1.313768278882945e+17, 1.313768278981382e+17, 1.313768279118883e+17, 1.313768279178257e+17, 1.313768279281382e+17, 1.313768279328257e+17, 1.31376827942982e+17, 1.313768279473571e+17, 1.313768279609508e+17, 1.313768279707945e+17, 1.31376827976732e+17, 1.313768279865757e+17, 1.313768279918883e+17, 1.313768280014195e+17, 1.313768280106382e+17, 1.31376828015482e+17, 1.313768280250132e+17, 1.313768280347008e+17, 1.313768280389196e+17, 1.31376828052982e+17, 1.313768280587631e+17, 1.31376828068607e+17, 1.313768280750132e+17, 1.313768280847007e+17, 1.31376828089857e+17, 1.31376828099857e+17, 1.313768281040758e+17, 1.313768281128257e+17, 1.313768281178258e+17, 1.313768281307945e+17, 1.313768281393883e+17, 1.313768281443882e+17, 1.313768281582945e+17, 1.31376828167982e+17, 1.313768281778257e+17, 1.313768281826694e+17, 1.313768281929819e+17, 1.313768282028257e+17, 1.313768282082945e+17, 1.31376828217982e+17, 1.313768282222007e+17, 1.313768282314195e+17, 1.313768282411071e+17, 1.313768282507945e+17, 1.313768282550132e+17, 1.313768282637633e+17, 1.31376828272357e+17, 1.313768282820444e+17, 1.31376828291732e+17, 1.313768282973569e+17, 1.313768283076695e+17, 1.313768283131382e+17, 1.313768283228257e+17, 1.313768283275133e+17, 1.313768283368882e+17, 1.313768283465757e+17, 1.313768283570445e+17, 1.313768283612632e+17, 1.313768283753257e+17, 1.313768283809508e+17, 1.313768283903258e+17, 1.313768283945445e+17, 1.313768284039195e+17, 1.313768284142321e+17, 1.313768284270445e+17, 1.313768284314195e+17, 1.313768284411071e+17, 1.313768284507945e+17, 1.313768284550134e+17, 1.313768284651695e+17, 1.313768284742319e+17, 1.313768284793883e+17, 1.313768284890757e+17, 1.313768284987633e+17, 1.31376828503607e+17, 1.313768285140758e+17, 1.313768285182945e+17, 1.313768285287633e+17, 1.31376828538607e+17, 1.313768285442319e+17, 1.313768285543882e+17, 1.31376828558607e+17, 1.313768285672008e+17, 1.313768285764195e+17, 1.31376828586732e+17, 1.313768285965757e+17, 1.313768286028257e+17, 1.313768286131383e+17, 1.313768286187633e+17, 1.31376828622982e+17, 1.31376828631732e+17, 1.313768286403258e+17, 1.313768286531383e+17, 1.313768286575132e+17, 1.313768286662632e+17, 1.31376828674857e+17, 1.313768286834509e+17, 1.313768286926696e+17, 1.31376828701732e+17, 1.313768287114195e+17, 1.313768287173569e+17, 1.313768287276695e+17, 1.313768287320445e+17, 1.313768287406382e+17, 1.31376828750482e+17, 1.313768287604819e+17, 1.313768287701695e+17, 1.313768287762632e+17, 1.31376828786107e+17, 1.313768287907945e+17, 1.313768288011069e+17, 1.313768288109508e+17, 1.31376828816732e+17, 1.313768288209508e+17, 1.313768288350132e+17, 1.313768288395446e+17, 1.313768288489194e+17, 1.313768288531383e+17, 1.31376828858607e+17, 1.313768288720444e+17, 1.31376828881732e+17, 1.313768288915757e+17, 1.313768288962633e+17, 1.313768289064196e+17, 1.313768289106383e+17, 1.31376828919232e+17, 1.313768289290757e+17, 1.313768289376695e+17, 1.313768289462633e+17, 1.313768289559507e+17, 1.313768289659508e+17, 1.313768289701696e+17, 1.313768289806383e+17, 1.313768289914195e+17, 1.313768290025133e+17, 1.313768290068882e+17, 1.313768290172008e+17, 1.313768290270445e+17, 1.313768290373569e+17, 1.313768290420445e+17, 1.313768290528257e+17, 1.313768290625133e+17, 1.313768290728257e+17, 1.313768290775132e+17, 1.313768290878257e+17, 1.313768290975132e+17, 1.313768291020445e+17, 1.313768291150132e+17, 1.31376829119232e+17, 1.313768291278258e+17, 1.313768291418883e+17, 1.313768291470445e+17, 1.313768291568882e+17, 1.313768291626694e+17, 1.31376829172357e+17, 1.313768291820444e+17, 1.313768291875132e+17, 1.31376829196107e+17, 1.313768292047008e+17, 1.313768292139195e+17, 1.313768292226694e+17, 1.313768292312632e+17, 1.313768292453258e+17, 1.313768292501695e+17, 1.313768292601695e+17, 1.31376829269857e+17, 1.313768292747008e+17, 1.313768292847007e+17, 1.313768292945445e+17, 1.31376829299232e+17, 1.313768293081382e+17, 1.31376829317982e+17, 1.313768293222007e+17, 1.313768293325133e+17, 1.313768293422008e+17, 1.313768293475132e+17, 1.313768293573571e+17, 1.313768293672008e+17, 1.313768293737633e+17, 1.31376829377982e+17, 1.313768293875133e+17, 1.313768293975132e+17, 1.313768294072008e+17, 1.313768294120445e+17, 1.31376829422982e+17, 1.313768294276695e+17, 1.313768294381382e+17, 1.31376829442357e+17, 1.313768294525133e+17, 1.313768294626694e+17, 1.313768294668882e+17, 1.313768294759507e+17, 1.313768294845444e+17, 1.313768294984507e+17, 1.313768295026694e+17, 1.31376829516107e+17, 1.313768295222007e+17, 1.313768295315758e+17, 1.313768295414195e+17, 1.313768295514195e+17, 1.313768295562632e+17, 1.31376829566107e+17, 1.313768295757946e+17, 1.313768295853257e+17, 1.313768295900133e+17, 1.31376829598607e+17, 1.313768296125133e+17, 1.313768296172008e+17, 1.313768296265757e+17, 1.313768296364195e+17, 1.313768296407945e+17, 1.31376829650482e+17, 1.313768296597009e+17, 1.313768296640758e+17, 1.313768296734508e+17, 1.31376829683607e+17, 1.313768296878258e+17, 1.313768297025133e+17, 1.313768297126696e+17, 1.313768297226694e+17, 1.313768297273571e+17, 1.313768297370445e+17, 1.31376829746732e+17, 1.313768297515758e+17, 1.313768297614195e+17, 1.313768297656383e+17, 1.313768297712632e+17, 1.313768297840756e+17, 1.313768297900133e+17, 1.313768298039195e+17, 1.31376829813607e+17, 1.313768298178257e+17, 1.313768298318883e+17, 1.313768298381382e+17, 1.31376829842357e+17, 1.313768298509508e+17, 1.31376829856732e+17, 1.313768298700133e+17, 1.313768298800132e+17, 1.313768298897007e+17, 1.313768298943882e+17, 1.313768299043882e+17, 1.313768299087633e+17, 1.313768299173571e+17, 1.313768299264196e+17, 1.313768299357944e+17, 1.313768299459507e+17, 1.313768299503258e+17, 1.313768299645445e+17, 1.31376829969232e+17, 1.313768299778257e+17, 1.313768299865757e+17, 1.313768299993883e+17, 1.313768300090757e+17, 1.313768300132946e+17, 1.313768300275132e+17, 1.313768300331382e+17, 1.31376830043607e+17, 1.313768300478258e+17, 1.313768300620444e+17, 1.313768300662633e+17, 1.313768300750132e+17, 1.313768300847007e+17, 1.31376830094857e+17, 1.313768300990757e+17, 1.313768301087633e+17, 1.313768301190757e+17, 1.313768301281382e+17, 1.31376830136732e+17, 1.313768301457946e+17, 1.313768301556383e+17, 1.31376830165482e+17, 1.313768301704819e+17, 1.313768301807945e+17, 1.313768301904819e+17, 1.31376830194857e+17, 1.313768302045445e+17, 1.313768302131383e+17, 1.31376830221732e+17, 1.31376830226732e+17, 1.313768302395444e+17, 1.313768302482945e+17, 1.313768302573569e+17, 1.31376830266732e+17, 1.313768302753257e+17, 1.313768302840756e+17, 1.313768302926696e+17, 1.313768303014195e+17, 1.31376830310482e+17, 1.313768303203258e+17, 1.313768303245445e+17, 1.313768303387633e+17, 1.313768303439195e+17, 1.313768303531382e+17, 1.31376830362982e+17, 1.31376830367982e+17, 1.313768303765757e+17, 1.313768303906383e+17, 1.31376830394857e+17, 1.313768304047008e+17, 1.313768304142321e+17, 1.31376830422982e+17, 1.31376830432357e+17, 1.313768304418883e+17, 1.313768304478257e+17, 1.313768304575132e+17, 1.313768304618883e+17, 1.313768304704819e+17, 1.313768304795444e+17, 1.313768304889196e+17, 1.313768304975132e+17, 1.313768305115757e+17, 1.313768305162633e+17, 1.313768305257944e+17, 1.313768305343882e+17, 1.313768305486071e+17, 1.313768305540758e+17, 1.313768305640756e+17, 1.313768305742319e+17, 1.313768305840758e+17, 1.31376830589232e+17, 1.313768305989196e+17, 1.313768306086071e+17, 1.31376830613607e+17, 1.313768306232945e+17, 1.31376830632982e+17, 1.313768306372008e+17, 1.313768306512632e+17, 1.31376830655482e+17, 1.313768306659507e+17, 1.313768306701695e+17, 1.313768306801695e+17, 1.313768306895446e+17, 1.313768306993883e+17, 1.313768307040758e+17, 1.313768307137633e+17, 1.313768307234509e+17, 1.313768307278258e+17, 1.313768307364196e+17, 1.313768307450132e+17, 1.31376830754857e+17, 1.313768307640758e+17, 1.313768307682945e+17, 1.313768307740758e+17, 1.313768307875132e+17, 1.313768307970445e+17, 1.313768308064195e+17, 1.313768308164196e+17, 1.313768308220445e+17, 1.313768308315758e+17, 1.313768308357946e+17, 1.31376830850482e+17, 1.313768308547008e+17, 1.313768308636069e+17, 1.313768308747008e+17, 1.313768308850132e+17, 1.313768308948571e+17, 1.313768308995444e+17, 1.31376830909232e+17, 1.313768309189194e+17, 1.313768309231382e+17, 1.31376830932982e+17, 1.313768309415758e+17, 1.313768309507945e+17, 1.313768309611071e+17, 1.313768309707945e+17, 1.31376830975482e+17, 1.31376830986732e+17, 1.313768309909508e+17, 1.313768310015757e+17, 1.313768310118883e+17, 1.313768310175133e+17, 1.313768310272008e+17, 1.313768310315757e+17, 1.313768310407945e+17, 1.313768310509508e+17, 1.313768310609507e+17, 1.31376831066107e+17, 1.313768310747008e+17, 1.313768310843884e+17, 1.313768310940758e+17, 1.313768311036069e+17, 1.313768311131383e+17, 1.313768311231383e+17, 1.313768311325133e+17, 1.313768311426696e+17, 1.31376831152357e+17, 1.31376831162357e+17, 1.313768311670445e+17, 1.313768311759507e+17, 1.313768311862633e+17, 1.313768311909508e+17, 1.313768312006382e+17, 1.313768312097007e+17, 1.313768312139195e+17, 1.313768312225133e+17, 1.313768312276695e+17, 1.313768312415758e+17, 1.313768312512632e+17, 1.313768312556383e+17, 1.313768312614195e+17, 1.313768312756383e+17, 1.313768312853258e+17, 1.313768312918883e+17, 1.313768313014195e+17, 1.313768313072008e+17, 1.313768313173569e+17, 1.313768313226694e+17, 1.313768313320444e+17, 1.31376831342357e+17, 1.313768313465757e+17, 1.313768313607945e+17, 1.313768313650132e+17, 1.313768313790757e+17, 1.313768313839195e+17, 1.313768313932945e+17, 1.313768313975132e+17, 1.313768314117321e+17, 1.313768314176695e+17, 1.313768314275133e+17, 1.313768314325133e+17, 1.313768314418883e+17, 1.313768314518883e+17, 1.313768314570445e+17, 1.313768314675132e+17, 1.313768314718883e+17, 1.313768314807945e+17, 1.31376831490482e+17, 1.31376831500482e+17, 1.313768315047008e+17, 1.313768315103258e+17, 1.313768315247008e+17, 1.313768315343882e+17, 1.31376831538607e+17, 1.313768315482944e+17, 1.313768315584507e+17, 1.313768315626696e+17, 1.313768315815757e+17, 1.313768315964196e+17, 1.313768316107944e+17, 1.313768316157946e+17, 1.313768316251695e+17, 1.313768316295444e+17, 1.31376831638607e+17, 1.313768316481382e+17, 1.313768316578258e+17, 1.313768316620445e+17, 1.313768316706382e+17, 1.313768316793883e+17, 1.313768316934508e+17, 1.313768316976695e+17, 1.31376831707982e+17, 1.313768317179821e+17, 1.313768317222008e+17, 1.313768317309508e+17, 1.313768317403258e+17, 1.31376831750482e+17, 1.313768317547007e+17, 1.313768317689196e+17, 1.313768317731383e+17, 1.313768317818883e+17, 1.313768317912632e+17, 1.313768318011071e+17, 1.31376831805482e+17, 1.313768318200133e+17, 1.313768318254821e+17, 1.313768318297007e+17, 1.31376831839232e+17, 1.313768318484507e+17, 1.313768318587633e+17, 1.313768318637633e+17, 1.313768318734508e+17, 1.31376831882982e+17, 1.313768318920444e+17, 1.313768319018883e+17, 1.313768319062633e+17, 1.31376831914857e+17, 1.313768319237632e+17, 1.313768319340758e+17, 1.313768319382944e+17, 1.31376831951732e+17, 1.313768319611069e+17, 1.313768319707945e+17, 1.313768319756383e+17, 1.313768319853257e+17, 1.313768319943882e+17, 1.313768320043882e+17, 1.313768320095444e+17, 1.31376832019232e+17, 1.313768320237632e+17, 1.313768320342319e+17, 1.313768320384507e+17, 1.313768320528257e+17, 1.313768320584508e+17, 1.31376832068607e+17, 1.313768320734508e+17, 1.31376832083607e+17, 1.313768320878258e+17, 1.313768320965757e+17, 1.31376832105482e+17, 1.313768321159508e+17, 1.313768321256383e+17, 1.313768321303258e+17, 1.313768321407945e+17, 1.31376832149857e+17, 1.31376832155482e+17, 1.313768321657944e+17, 1.313768321700133e+17, 1.313768321790758e+17, 1.31376832188607e+17, 1.313768321984508e+17, 1.313768322031382e+17, 1.313768322137633e+17, 1.313768322179821e+17, 1.31376832226732e+17, 1.313768322315757e+17, 1.313768322443882e+17, 1.313768322534508e+17, 1.313768322628257e+17, 1.313768322731383e+17, 1.313768322773571e+17, 1.31376832286732e+17, 1.313768322968883e+17, 1.313768323065757e+17, 1.313768323114195e+17, 1.313768323212634e+17, 1.313768323311069e+17, 1.313768323409508e+17, 1.313768323465757e+17, 1.313768323557946e+17, 1.313768323603258e+17, 1.313768323695444e+17, 1.313768323795444e+17, 1.313768323890757e+17, 1.313768323940758e+17, 1.31376832403607e+17, 1.313768324128257e+17, 1.313768324228257e+17, 1.313768324322007e+17, 1.313768324364195e+17, 1.313768324451695e+17, 1.313768324545444e+17, 1.313768324650132e+17, 1.313768324750132e+17, 1.313768324847008e+17, 1.313768324906383e+17, 1.31376832500482e+17, 1.313768325056383e+17, 1.313768325164196e+17, 1.313768325206382e+17, 1.31376832526107e+17, 1.313768325389196e+17, 1.313768325476695e+17, 1.313768325562633e+17, 1.313768325651694e+17, 1.313768325740758e+17, 1.313768325828257e+17, 1.313768325918883e+17, 1.313768326018883e+17, 1.31376832606107e+17, 1.31376832616732e+17, 1.313768326259507e+17, 1.313768326306382e+17, 1.313768326411069e+17, 1.313768326509508e+17, 1.313768326551694e+17, 1.313768326643882e+17, 1.313768326737633e+17, 1.313768326839196e+17, 1.313768326881382e+17, 1.313768326968883e+17, 1.313768327059507e+17, 1.313768327162633e+17, 1.313768327253257e+17, 1.313768327295446e+17, 1.313768327382944e+17, 1.313768327468882e+17, 1.313768327607945e+17, 1.313768327706382e+17, 1.313768327757946e+17, 1.313768327856383e+17, 1.313768327953257e+17, 1.313768328007945e+17},
			             {1.313768170672008e+17, 1.313768171156383e+17},
			             {1.313768117743882e+17, 1.313768118395444e+17},
			             {1.313768119626694e+17, 1.313768119870445e+17},
			             {1.31376812029857e+17, 1.313768120401696e+17},
			             {1.313768120743882e+17, 1.313768120928257e+17},
			             {1.313768122351695e+17, 1.31376812289232e+17},
			             {1.313768126386071e+17, 1.313768126514195e+17},
			             {1.313768128932945e+17, 1.313768129303258e+17},
			             {1.313768184926696e+17, 1.313768185526696e+17},
			             {1.313768190501695e+17, 1.31376819063607e+17},
			             {1.31376825916732e+17, 1.31376825996107e+17},
			             {1.313768278647008e+17, 1.313768279118883e+17},
			             {1.313768289914195e+17, 1.313768291020445e+17},
			             {1.31376829317982e+17, 1.313768293325133e+17},
			             {1.313768296172008e+17, 1.313768296265757e+17, 1.313768296364195e+17, 1.313768296407945e+17, 1.31376829650482e+17, 1.313768296597009e+17, 1.313768296640758e+17, 1.313768296734508e+17, 1.31376829683607e+17, 1.313768296878258e+17, 1.313768297025133e+17, 1.313768297126696e+17, 1.313768297226694e+17, 1.313768297273571e+17, 1.313768297370445e+17, 1.31376829746732e+17, 1.313768297515758e+17, 1.313768297614195e+17, 1.313768297656383e+17, 1.313768297712632e+17, 1.313768297840756e+17, 1.313768298381382e+17},
			             {1.31376828167982e+17},
			             {1.313768279707945e+17, 1.313768280106382e+17},
			             {1.313768328007945e+17},
			             {1.313768256725133e+17, 1.31376825712982e+17},
			             {1.313768212506383e+17, 1.313768212548571e+17},
			             {1.313768327382944e+17, 1.313768327706382e+17};
			mask_depths = {{15.0, 15.0, 71.0, 71.0}, {15.0, 71.1}, {15.0, 71.2}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.2}, {15.0, 71.2}, {15.0, 71.2}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.7}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.4}, {15.0, 72.5}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.9}, {15.0, 72.8}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.3}, {15.0, 72.1}, {15.0, 72.0}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.3}, {15.0, 71.2}, {15.0, 71.1}, {15.0, 70.9}, {15.0, 70.9}, {15.0, 70.8}, {15.0, 70.8}, {15.0, 70.9}, {15.0, 71.2}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 71.9}, {15.0, 71.6}, {15.0, 71.4}, {15.0, 71.2}, {15.0, 71.1}, {15.0, 71.2}, {15.0, 71.4}, {15.0, 71.8}, {15.0, 72.0}, {15.0, 72.1}, {15.0, 72.4}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.5}, {15.0, 72.4}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.6}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.1}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 71.7}, {15.0, 71.6}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.7}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 71.7}, {15.0, 71.5}, {15.0, 71.2}, {15.0, 71.1}, {15.0, 71.0}, {15.0, 70.9}, {15.0, 71.1}, {15.0, 71.4}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 72.2}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 71.8}, {15.0, 71.5}, {15.0, 71.2}, {15.0, 71.1}, {15.0, 71.2}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.2}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 71.1}, {15.0, 71.0}, {15.0, 70.9}, {15.0, 70.7}, {15.0, 70.6}, {15.0, 70.4}, {15.0, 70.3}, {15.0, 70.4}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.6}, {15.0, 70.6}, {15.0, 70.4}, {15.0, 70.4}, {15.0, 70.5}, {15.0, 70.4}, {15.0, 70.4}, {15.0, 70.3}, {15.0, 70.2}, {15.0, 70.3}, {15.0, 70.5}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.6}, {15.0, 70.5}, {15.0, 70.4}, {15.0, 70.4}, {15.0, 70.4}, {15.0, 70.4}, {15.0, 70.4}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.6}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.9}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 70.9}, {15.0, 70.9}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 71.2}, {15.0, 71.2}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.1}, {15.0, 71.1}, {15.0, 71.1}, {15.0, 71.2}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.7}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.7}, {15.0, 71.9}, {15.0, 71.9}, {15.0, 71.9}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.7}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 72.0}, {15.0, 72.2}, {15.0, 72.4}, {15.0, 72.5}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.7}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.7}, {15.0, 72.6}, {15.0, 72.7}, {15.0, 72.6}, {15.0, 72.7}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.3}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.7}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 73.1}, {15.0, 73.1}, {15.0, 73.4}, {15.0, 73.7}, {15.0, 73.9}, {15.0, 73.9}, {15.0, 73.9}, {15.0, 73.9}, {15.0, 73.8}, {15.0, 73.8}, {15.0, 73.7}, {15.0, 73.6}, {15.0, 73.6}, {15.0, 73.7}, {15.0, 73.7}, {15.0, 73.5}, {15.0, 73.4}, {15.0, 73.4}, {15.0, 72.8}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.8}, {15.0, 72.9}, {15.0, 73.1}, {15.0, 73.1}, {15.0, 73.1}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.1}, {15.0, 72.8}, {15.0, 72.6}, {15.0, 72.0}, {15.0, 71.9}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.1}, {15.0, 71.2}, {15.0, 71.2}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.2}, {15.0, 71.0}, {15.0, 70.8}, {15.0, 70.7}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.6}, {15.0, 70.6}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.8}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.5}, {15.0, 70.5}, {15.0, 70.5}, {15.0, 70.4}, {15.0, 70.6}, {15.0, 70.9}, {15.0, 71.1}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 72.0}, {15.0, 72.6}, {15.0, 72.1}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 71.9}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.1}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.5}, {15.0, 72.8}, {15.0, 72.9}, {15.0, 73.0}, {15.0, 73.0}, {15.0, 72.9}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.9}, {15.0, 73.0}, {15.0, 73.1}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.1}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.9}, {15.0, 73.1}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.1}, {15.0, 72.9}, {15.0, 72.8}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.7}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 73.0}, {15.0, 73.0}, {15.0, 73.0}, {15.0, 73.0}, {15.0, 72.7}, {15.0, 72.8}, {15.0, 72.9}, {15.0, 72.9}, {15.0, 73.1}, {15.0, 73.2}, {15.0, 73.3}, {15.0, 73.4}, {15.0, 73.7}, {15.0, 73.9}, {15.0, 73.9}, {15.0, 73.6}, {15.0, 73.6}, {15.0, 73.3}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.3}, {15.0, 73.6}, {15.0, 73.6}, {15.0, 73.7}, {15.0, 73.8}, {15.0, 73.8}, {15.0, 73.9}, {15.0, 73.8}, {15.0, 73.9}, {15.0, 73.8}, {15.0, 73.9}, {15.0, 74.0}, {15.0, 74.0}, {15.0, 74.2}, {15.0, 74.2}, {15.0, 74.2}, {15.0, 74.1}, {15.0, 73.7}, {15.0, 73.6}, {15.0, 73.3}, {15.0, 73.3}, {15.0, 73.2}, {15.0, 73.1}, {15.0, 73.0}, {15.0, 73.0}, {15.0, 72.9}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.7}, {15.0, 72.6}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.5}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.5}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.9}, {15.0, 73.1}, {15.0, 73.1}, {15.0, 73.2}, {15.0, 73.4}, {15.0, 73.5}, {15.0, 73.6}, {15.0, 73.6}, {15.0, 73.7}, {15.0, 73.8}, {15.0, 73.8}, {15.0, 73.9}, {15.0, 73.9}, {15.0, 73.9}, {15.0, 73.7}, {15.0, 73.6}, {15.0, 73.5}, {15.0, 73.5}, {15.0, 73.5}, {15.0, 73.6}, {15.0, 73.5}, {15.0, 73.4}, {15.0, 73.3}, {15.0, 73.2}, {15.0, 73.0}, {15.0, 72.8}, {15.0, 72.8}, {15.0, 72.9}, {15.0, 72.9}, {15.0, 72.9}, {15.0, 73.0}, {15.0, 73.0}, {15.0, 72.9}, {15.0, 72.7}, {15.0, 72.6}, {15.0, 72.5}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.8}, {15.0, 72.7}, {15.0, 72.5}, {15.0, 72.4}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.8}, {15.0, 73.0}, {15.0, 73.2}, {15.0, 73.3}, {15.0, 73.3}, {15.0, 73.2}, {15.0, 73.1}, {15.0, 73.0}, {15.0, 73.0}, {15.0, 73.1}, {15.0, 73.5}, {15.0, 73.6}, {15.0, 73.9}, {15.0, 74.0}, {15.0, 74.1}, {15.0, 74.2}, {15.0, 74.1}, {15.0, 74.1}, {15.0, 73.9}, {15.0, 73.9}, {15.0, 74.0}, {15.0, 74.0}, {15.0, 73.9}, {15.0, 73.8}, {15.0, 73.7}, {15.0, 73.5}, {15.0, 73.4}, {15.0, 73.4}, {15.0, 73.4}, {15.0, 73.5}, {15.0, 73.5}, {15.0, 73.5}, {15.0, 73.5}, {15.0, 73.6}, {15.0, 73.5}, {15.0, 73.7}, {15.0, 73.8}, {15.0, 73.8}, {15.0, 73.8}, {15.0, 73.8}, {15.0, 73.8}, {15.0, 73.8}, {15.0, 73.6}, {15.0, 73.6}, {15.0, 73.6}, {15.0, 73.7}, {15.0, 73.7}, {15.0, 73.7}, {15.0, 73.6}, {15.0, 73.4}, {15.0, 73.3}, {15.0, 73.0}, {15.0, 72.7}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 73.0}, {15.0, 73.3}, {15.0, 73.3}, {15.0, 73.4}, {15.0, 73.3}, {15.0, 73.3}, {15.0, 73.3}, {15.0, 73.2}, {15.0, 73.3}, {15.0, 73.6}, {15.0, 74.1}, {15.0, 74.2}, {15.0, 74.4}, {15.0, 74.6}, {15.0, 74.7}, {15.0, 74.7}, {15.0, 74.7}, {15.0, 74.6}, {15.0, 74.5}, {15.0, 74.7}, {15.0, 74.7}, {15.0, 74.8}, {15.0, 74.9}, {15.0, 75.0}, {15.0, 75.0}, {15.0, 74.8}, {15.0, 74.5}, {15.0, 74.1}, {15.0, 73.9}, {15.0, 73.7}, {15.0, 73.6}, {15.0, 73.5}, {15.0, 73.3}, {15.0, 73.1}, {15.0, 72.7}, {15.0, 72.5}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.1}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 71.9}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.3}, {15.0, 71.2}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 71.1}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.2}, {15.0, 71.5}, {15.0, 71.7}, {15.0, 71.9}, {15.0, 72.0}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 71.9}, {15.0, 72.1}, {15.0, 72.5}, {15.0, 72.8}, {15.0, 73.0}, {15.0, 73.1}, {15.0, 73.6}, {15.0, 74.0}, {15.0, 74.2}, {15.0, 74.1}, {15.0, 74.1}, {15.0, 74.1}, {15.0, 74.1}, {15.0, 74.2}, {15.0, 74.1}, {15.0, 74.0}, {15.0, 73.9}, {15.0, 73.6}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 72.9}, {15.0, 72.7}, {15.0, 72.5}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.2}, {15.0, 71.2}, {15.0, 71.7}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 72.0}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 71.9}, {15.0, 72.0}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 71.9}, {15.0, 71.9}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.7}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.3}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 71.9}, {15.0, 72.0}, {15.0, 72.1}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.0}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.4}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.0}, {15.0, 72.0}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 72.0}, {15.0, 72.1}, {15.0, 72.1}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 72.0}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.7}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.0}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.8}, {15.0, 71.3}, {15.0, 71.3}, {15.0, 71.5}, {15.0, 71.7}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.5}, {15.0, 72.8}, {15.0, 73.0}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.2}, {15.0, 73.1}, {15.0, 72.9}, {15.0, 72.7}, {15.0, 72.6}, {15.0, 72.5}, {15.0, 72.4}, {15.0, 72.2}, {15.0, 71.9}, {15.0, 71.6}, {15.0, 71.3}, {15.0, 71.1}, {15.0, 70.8}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.6}, {15.0, 70.5}, {15.0, 70.5}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.2}, {15.0, 70.2}, {15.0, 70.3}, {15.0, 70.4}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.0}, {15.0, 69.9}, {15.0, 69.8}, {15.0, 69.5}, {15.0, 69.6}, {15.0, 69.6}, {15.0, 69.9}, {15.0, 70.0}, {15.0, 70.2}, {15.0, 70.2}, {15.0, 70.3}, {15.0, 70.2}, {15.0, 70.2}, {15.0, 70.1}, {15.0, 70.1}, {15.0, 70.1}, {15.0, 70.1}, {15.0, 70.1}, {15.0, 70.2}, {15.0, 70.2}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.2}, {15.0, 70.0}, {15.0, 69.9}, {15.0, 69.7}, {15.0, 69.7}, {15.0, 69.8}, {15.0, 70.0}, {15.0, 70.4}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.7}, {15.0, 70.8}, {15.0, 70.8}, {15.0, 70.8}, {15.0, 70.8}, {15.0, 70.9}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 71.1}, {15.0, 71.1}, {15.0, 71.1}, {15.0, 71.0}, {15.0, 70.9}, {15.0, 70.8}, {15.0, 70.8}, {15.0, 70.6}, {15.0, 70.7}, {15.0, 70.6}, {15.0, 70.6}, {15.0, 70.5}, {15.0, 70.5}, {15.0, 70.4}, {15.0, 70.4}, {15.0, 70.3}, {15.0, 70.2}, {15.0, 70.1}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 70.2}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.1}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 70.1}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.3}, {15.0, 70.2}, {15.0, 70.1}, {15.0, 70.1}, {15.0, 70.1}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 69.9}, {15.0, 69.8}, {15.0, 69.8}, {15.0, 70.0}, {15.0, 70.4}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.8}, {15.0, 71.0}, {15.0, 71.1}, {15.0, 71.1}, {15.0, 71.1}, {15.0, 71.4}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 71.9}, {15.0, 72.1}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.2}, {15.0, 72.0}, {15.0, 71.9}, {15.0, 71.8}, {15.0, 71.8}, {15.0, 71.5}, {15.0, 71.5}, {15.0, 71.2}, {15.0, 70.9}, {15.0, 70.7}, {15.0, 70.5}, {15.0, 70.4}, {15.0, 70.1}, {15.0, 70.1}, {15.0, 69.9}, {15.0, 69.8}, {15.0, 69.6}, {15.0, 69.5}, {15.0, 69.4}, {15.0, 69.4}, {15.0, 69.3}, {15.0, 69.4}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.2}, {15.0, 69.1}, {15.0, 69.0}, {15.0, 68.8}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.8}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.4}, {15.0, 69.5}, {15.0, 69.5}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.4}, {15.0, 69.6}, {15.0, 69.8}, {15.0, 69.8}, {15.0, 69.8}, {15.0, 69.8}, {15.0, 69.6}, {15.0, 69.5}, {15.0, 69.3}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.5}, {15.0, 69.7}, {15.0, 70.0}, {15.0, 70.1}, {15.0, 70.3}, {15.0, 70.4}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.5}, {15.0, 70.6}, {15.0, 70.6}, {15.0, 70.6}, {15.0, 70.8}, {15.0, 70.7}, {15.0, 70.6}, {15.0, 70.4}, {15.0, 70.1}, {15.0, 70.0}, {15.0, 69.8}, {15.0, 69.7}, {15.0, 69.6}, {15.0, 69.7}, {15.0, 69.7}, {15.0, 69.6}, {15.0, 69.5}, {15.0, 69.4}, {15.0, 69.2}, {15.0, 69.0}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.7}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 69.4}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.4}, {15.0, 69.4}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.2}, {15.0, 69.1}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 69.1}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.0}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.6}, {15.0, 69.7}, {15.0, 69.7}, {15.0, 69.7}, {15.0, 69.8}, {15.0, 69.8}, {15.0, 69.9}, {15.0, 69.9}, {15.0, 70.1}, {15.0, 70.3}, {15.0, 70.4}, {15.0, 70.4}, {15.0, 70.2}, {15.0, 70.2}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 69.8}, {15.0, 69.8}, {15.0, 70.3}, {15.0, 70.5}, {15.0, 70.8}, {15.0, 71.2}, {15.0, 71.4}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.3}, {15.0, 71.2}, {15.0, 71.1}, {15.0, 71.1}, {15.0, 71.0}, {15.0, 70.8}, {15.0, 70.7}, {15.0, 70.4}, {15.0, 70.0}, {15.0, 69.8}, {15.0, 69.5}, {15.0, 69.3}, {15.0, 69.2}, {15.0, 69.1}, {15.0, 69.1}, {15.0, 68.9}, {15.0, 68.6}, {15.0, 68.3}, {15.0, 68.1}, {15.0, 67.8}, {15.0, 67.4}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 68.1}, {15.0, 68.2}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.6}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.1}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.4}, {15.0, 69.4}, {15.0, 69.4}, {15.0, 69.3}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 68.8}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.5}, {15.0, 68.3}, {15.0, 68.2}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.1}, {15.0, 67.0}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 67.0}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.1}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 67.1}, {15.0, 67.5}, {15.0, 67.6}, {15.0, 68.1}, {15.0, 68.4}, {15.0, 68.5}, {15.0, 68.7}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 68.7}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.2}, {15.0, 68.2}, {15.0, 68.1}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.2}, {15.0, 67.1}, {15.0, 67.0}, {15.0, 66.8}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.4}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.3}, {15.0, 66.6}, {15.0, 66.9}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.0}, {15.0, 66.8}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 67.0}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 67.9}, {15.0, 68.2}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.0}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.4}, {15.0, 66.4}, {15.0, 66.3}, {15.0, 66.6}, {15.0, 66.9}, {15.0, 67.1}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 68.0}, {15.0, 68.2}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.2}, {15.0, 68.1}, {15.0, 67.7}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.5}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.4}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.3}, {15.0, 66.4}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.4}, {15.0, 66.4}, {15.0, 66.4}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.2}, {15.0, 66.2}, {15.0, 66.4}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.1}, {15.0, 67.0}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.6}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 67.9}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 67.9}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 68.0}, {15.0, 68.2}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.5}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.2}, {15.0, 68.5}, {15.0, 68.7}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.1}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.1}, {15.0, 69.2}, {15.0, 69.1}, {15.0, 69.1}, {15.0, 69.0}, {15.0, 68.9}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.5}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.2}, {15.0, 68.0}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.7}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 68.3}, {15.0, 68.2}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 68.1}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 69.1}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.2}, {15.0, 69.1}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.4}, {15.0, 69.5}, {15.0, 69.5}, {15.0, 69.5}, {15.0, 69.5}, {15.0, 69.4}, {15.0, 69.0}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 68.8}, {15.0, 68.7}, {15.0, 68.2}, {15.0, 67.8}, {15.0, 67.6}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 68.4}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.0}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.2}, {15.0, 68.2}, {15.0, 68.2}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.2}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.2}, {15.0, 68.2}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.1}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.5}, {15.0, 67.6}, {15.0, 67.8}, {15.0, 70.7}, {15.0, 68.4}, {15.0, 68.6}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 68.9}, {15.0, 68.8}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.2}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.7}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.2}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 67.0}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.7}, {15.0, 68.1}, {15.0, 68.4}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.4}, {15.0, 68.2}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.1}, {15.0, 66.9}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 68.5}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.7}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.3}, {15.0, 68.2}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 67.9}, {15.0, 67.7}, {15.0, 67.5}, {15.0, 67.3}, {15.0, 67.0}, {15.0, 66.9}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.8}, {15.0, 67.0}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.6}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.1}, {15.0, 67.0}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.0}, {15.0, 66.8}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.4}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.1}, {15.0, 66.8}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.2}, {15.0, 66.3}, {15.0, 66.5}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.7}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.2}, {15.0, 67.5}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.7}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.0}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.4}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.4}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.4}, {15.0, 66.4}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.2}, {15.0, 66.1}, {15.0, 66.2}, {15.0, 66.4}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.1}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 67.0}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.2}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.2}, {15.0, 66.2}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.2}, {15.0, 66.2}, {15.0, 66.0}, {15.0, 65.9}, {15.0, 65.8}, {15.0, 65.7}, {15.0, 65.7}, {15.0, 65.8}, {15.0, 65.9}, {15.0, 66.1}, {15.0, 66.2}, {15.0, 66.3}, {15.0, 66.4}, {15.0, 66.2}, {15.0, 66.1}, {15.0, 65.9}, {15.0, 65.8}, {15.0, 65.7}, {15.0, 65.7}, {15.0, 66.0}, {15.0, 66.1}, {15.0, 66.4}, {15.0, 66.7}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.2}, {15.0, 68.2}, {15.0, 68.5}, {15.0, 68.9}, {15.5, 68.9}, {15.5, 69.2}, {15.5, 69.3}, {15.3, 69.3}, {15.2, 69.2}, {15.0, 69.1}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 68.8}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.4}, {15.0, 67.8}, {15.0, 67.6}, {15.0, 67.2}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.6}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.2}, {15.0, 66.1}, {15.0, 66.1}, {15.0, 66.1}, {15.0, 65.9}, {15.0, 65.7}, {15.0, 65.7}, {15.0, 65.5}, {15.0, 65.6}, {15.0, 65.7}, {15.0, 65.9}, {15.0, 66.0}, {15.0, 66.1}, {15.0, 66.2}, {15.0, 66.2}, {15.0, 66.2}, {15.0, 66.0}, {15.0, 65.9}, {15.0, 65.8}, {15.0, 65.7}, {15.0, 65.8}, {15.0, 65.9}, {15.0, 66.0}, {15.0, 66.2}, {15.0, 66.2}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.5}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.3}, {15.0, 66.5}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 67.0}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.0}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.5}, {15.0, 66.5}, {15.0, 66.4}, {15.0, 66.5}, {15.0, 66.6}, {15.0, 66.7}, {15.0, 66.7}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.9}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.4}, {15.0, 67.3}, {15.0, 67.1}, {15.0, 67.1}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.5}, {15.0, 67.6}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.5}, {15.0, 68.2}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.5}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.1}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.1}, {15.0, 69.1}, {15.0, 69.0}, {15.0, 68.9}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.5}, {15.0, 68.3}, {15.0, 68.2}, {15.0, 68.1}, {15.0, 68.1}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.6}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.2}, {15.0, 67.3}, {15.0, 67.2}, {15.0, 67.1}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 66.9}, {15.0, 67.2}, {15.0, 67.4}, {15.0, 67.5}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.7}, {15.0, 67.8}, {15.0, 67.7}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.6}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 67.8}, {15.0, 67.9}, {15.0, 67.9}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.0}, {15.0, 68.1}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.5}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 69.1}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.2}, {15.0, 69.0}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.5}, {15.0, 69.6}, {15.0, 69.7}, {15.0, 69.6}, {15.0, 69.5}, {15.0, 69.2}, {15.0, 69.1}, {15.0, 69.0}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.3}, {15.0, 69.4}, {15.0, 69.3}, {15.0, 69.1}, {15.0, 68.9}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.6}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.2}, {15.0, 68.3}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 68.8}, {15.0, 68.9}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 68.8}, {15.0, 68.8}, {15.0, 68.6}, {15.0, 68.7}, {15.0, 68.7}, {15.0, 69.0}, {15.0, 69.0}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.4}, {15.0, 69.5}, {15.0, 69.7}, {15.0, 69.8}, {15.0, 69.9}, {15.0, 70.0}, {15.0, 69.9}, {15.0, 69.9}, {15.0, 69.9}, {15.0, 69.8}, {15.0, 69.9}, {15.0, 70.6}, {15.0, 70.8}, {15.0, 70.9}, {17.1, 71.3}, {17.3, 71.8}, {17.7, 71.9}, {17.2, 72.3}, {16.0, 72.3}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.3}, {15.0, 72.1}, {15.0, 71.9}, {15.0, 71.5}, {15.0, 71.2}, {15.0, 70.9}, {15.0, 70.8}, {15.0, 70.5}, {15.0, 70.3}, {15.0, 69.9}, {15.0, 69.7}, {15.0, 69.5}, {15.0, 69.2}, {15.0, 69.1}, {15.0, 68.9}, {15.0, 68.7}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.5}, {15.0, 68.4}, {15.0, 68.4}, {15.0, 68.3}, {15.0, 68.4}, {15.0, 68.6}, {15.0, 68.9}, {15.0, 69.0}, {15.0, 69.2}, {15.0, 69.3}, {15.0, 69.5}, {15.0, 69.6}, {15.0, 69.6}, {15.0, 69.8}, {15.0, 69.8}, {15.0, 69.9}, {15.0, 69.8}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 69.9}, {15.0, 69.9}, {15.0, 69.8}, {15.0, 69.8}, {15.0, 69.9}, {15.0, 70.1}, {15.0, 70.1}, {15.0, 69.9}, {15.0, 70.1}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 70.0}, {15.0, 69.9}, {15.0, 70.1}, {15.0, 70.4}, {15.0, 70.6}, {15.0, 70.7}, {15.0, 70.8}, {15.0, 70.9}, {15.0, 70.9}, {15.0, 70.9}, {15.0, 70.8}, {15.0, 70.8}, {15.0, 71.0}, {15.0, 71.2}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 71.3}, {15.0, 71.5}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.6}, {15.0, 71.5}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.3}, {15.0, 71.2}, {15.0, 71.1}, {15.0, 71.2}, {15.0, 71.2}, {15.0, 71.1}, {15.0, 71.1}, {15.0, 71.0}, {15.0, 70.9}, {15.0, 70.8}, {15.0, 70.7}, {15.0, 70.7}, {15.0, 70.6}, {15.0, 70.7}, {15.0, 70.9}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 71.0}, {15.0, 70.9}, {15.0, 70.8}, {15.0, 70.8}, {15.0, 70.8}, {15.0, 70.9}, {15.0, 71.2}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.4}, {15.0, 71.5}, {15.0, 71.8}, {15.0, 71.9}, {15.0, 72.2}, {15.0, 72.3}, {15.0, 72.4}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.5}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.6}, {15.0, 72.7}, {15.0, 72.7}, {15.0, 72.6}, {15.0, 72.4}, {15.0, 72.4}, {15.0, 72.2}, {15.0, 72.1}, {15.0, 72.2}, {15.0, 72.5}, {15.0, 72.7}, {15.0, 72.4}, {15.0, 72.1}, {15.0, 15.0, 72.9, 72.9}}, {{21.2, 34.6}, {21.2, 34.6}}, {{20.7, 34.5}, {20.7, 34.5}}, {{19.9, 24.9}, {19.9, 24.9}}, {{24.3, 31.2}, {24.3, 31.2}}, {{19.2, 25.9}, {19.2, 25.9}}, {{17.3, 31.7}, {17.3, 31.7}}, {{18.8, 24.7}, {18.8, 24.7}}, {{18.6, 34.7}, {18.6, 34.7}}, {{27.2, 35.8}, {27.2, 35.8}}, {{27.1, 34.7}, {27.1, 34.7}}, {{35.5, 46.6}, {35.5, 46.6}}, {{25.9, 38.8}, {25.9, 38.8}}, {{28.9, 43.8}, {28.9, 43.8}}, {{33.6, 37.8}, {33.6, 37.8}}, {{37.8, 40.6, 40.8}, {36.3, 37.7, 40.5}, {36.0, 36.2}, {35.6, 35.9, 40.7, 40.9}, {35.1, 35.5, 41.0, 41.3}, {34.5, 35.0, 41.4, 41.5}, {33.9, 34.4}, {33.3, 33.8, 41.7, 42.2}, {32.8, 33.2, 42.3, 42.4}, {32.2, 32.7, 42.5, 43.3}, {43.4, 43.5}, {43.6}, {31.8, 31.9}, {31.6, 31.7}, {31.1, 31.5}, {30.7, 31.0}, {30.4, 30.6}, {30.0, 30.3}, {29.6, 29.9}, {28.8, 28.9, 29.5}, {29.0}, {29.0, 43.6}}, {{2.4, 2.4, 2.8, 2.8}}, {{63.1, 66.3}, {63.1, 66.3}}, {{3.9, 3.9, 4.1, 4.1}}, {{64.3, 67.7}, {64.3, 67.7}}, {{20.2, 22.5}, {20.2, 22.5}}, {{38.6, 45.2}, {38.6, 45.2}};
		}
	}
}
