netcdf mask {
	:date_created = "20200811T114628";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200811T114628";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 26;
			channels = 4;
			categories = 104;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  39.8, 39.9, 39.2, 39.1, 36.9, 38.9, 39.9, 40.2, 38.4, 37.6, 37.4, 37.4, 37.4, 37.5, 36.3, 36.4, 37.2, 37.0, 37.6, 36.5, 36.8, 30.0, 35.9, 21.9, 41.8, 42.3;
			max_depth =  42.9, 41.6, 41.0, 40.4, 40.2, 40.0, 40.9, 41.0, 39.6, 38.7, 38.5, 38.5, 38.5, 38.5, 37.7, 38.1, 38.0, 38.0, 38.6, 38.3, 38.8, 36.1, 38.8, 31.8, 44.9, 45.6;
			start_time = 129799100934102016, 129799101572695808, 129799101677070720, 129799101701133184, 129799101765352064, 129799101797539456, 129799101825664512, 129799101837695744, 129799101966289536, 129799101978320768, 129799102150977024, 129799102175039488, 129799102215195776, 129799102243320832, 129799102476289536, 129799102492383232, 129799102516445696, 129799102536445696, 129799102596758272, 129799102693164416, 129799102809570816, 129799102905976960, 129799102938164480, 129799117242851968, 129799106066445824, 129799106295352064;
			end_time = 129799100970195712, 129799101588789504, 129799101697070720, 129799101713164544, 129799101789570816, 129799101805664512, 129799101833633152, 129799101845820672, 129799101974258304, 129799101990352000, 129799102158945792, 129799102179102080, 129799102223320832, 129799102247383168, 129799102484258176, 129799102512383232, 129799102528476928, 129799102548477056, 129799102608789504, 129799102713164544, 129799102845664512, 129799102922070784, 129799102950195712, 129799117295195776, 129799106094570752, 129799106335664512;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21","Layer22","Layer23","Layer24","Layer25","Layer26";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "200", "333";
			region_channels = 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15;
			mask_times = {1.29799100934102e+17, 1.297991009420708e+17, 1.297991009461332e+17, 1.297991009501957e+17, 1.297991009542583e+17, 1.297991009701957e+17},
			             {1.297991015726958e+17, 1.29799101584727e+17, 1.297991015887895e+17},
			             {1.297991016770707e+17, 1.297991016970707e+17},
			             {1.297991017011332e+17, 1.297991017131645e+17},
			             {1.297991017653521e+17, 1.297991017694145e+17, 1.297991017775396e+17, 1.297991017855082e+17, 1.297991017895708e+17},
			             {1.297991017975395e+17, 1.297991018056645e+17},
			             {1.297991018256645e+17, 1.297991018336332e+17},
			             {1.297991018376957e+17, 1.297991018458207e+17},
			             {1.297991019662895e+17, 1.297991019742583e+17},
			             {1.297991019783208e+17, 1.29799101990352e+17},
			             {1.29799102150977e+17, 1.297991021589458e+17},
			             {1.297991021750395e+17, 1.297991021791021e+17},
			             {1.297991022151958e+17, 1.297991022233208e+17},
			             {1.297991022433208e+17, 1.297991022473832e+17},
			             {1.297991024762895e+17, 1.297991024842582e+17},
			             {1.297991024923832e+17, 1.297991025044145e+17, 1.297991025083208e+17, 1.297991025123832e+17},
			             {1.297991025164457e+17, 1.29799102520352e+17, 1.297991025244145e+17, 1.297991025284769e+17},
			             {1.297991025364457e+17, 1.297991025405083e+17, 1.297991025445708e+17, 1.297991025484771e+17},
			             {1.297991025967583e+17, 1.297991026008207e+17, 1.297991026087895e+17},
			             {1.297991026931644e+17, 1.297991027131645e+17},
			             {1.297991028095708e+17, 1.297991028256645e+17, 1.297991028295708e+17, 1.297991028376957e+17, 1.297991028456645e+17},
			             {1.29799102905977e+17, 1.297991029220708e+17},
			             {1.297991029381645e+17, 1.297991029461332e+17, 1.297991029501957e+17},
			             {1.29799117242852e+17, 1.297991172951958e+17},
			             {1.297991060664458e+17, 1.297991060705083e+17, 1.297991060786333e+17, 1.29799106086602e+17, 1.297991060945708e+17},
			             {1.297991062953521e+17, 1.29799106303477e+17, 1.297991063075396e+17, 1.297991063155084e+17, 1.297991063195707e+17, 1.29799106323477e+17, 1.297991063275396e+17, 1.297991063316019e+17, 1.297991063356645e+17};
			mask_depths = {{39.8, 42.9}, {42.9}, {42.8}, {42.8}, {42.7}, {39.8, 42.7}}, {{39.9, 41.6}, {41.6}, {39.9, 41.5}}, {{39.2, 41.0}, {39.2, 41.0}}, {{39.1, 40.4}, {39.1, 40.4}}, {{36.9, 40.2}, {40.2}, {40.0}, {40.0}, {36.9, 40.1}}, {{38.9, 40.0}, {38.9, 40.0}}, {{39.9, 40.7}, {39.9, 40.9}}, {{40.2, 41.0}, {40.2, 41.0}}, {{38.4, 39.6}, {38.4, 39.6}}, {{37.6, 38.7}, {37.6, 38.7}}, {{37.4, 38.5}, {37.4, 38.5}}, {{37.4, 38.5}, {37.4, 38.5}}, {{37.4, 38.5}, {37.4, 38.5}}, {{37.5, 38.5}, {37.5, 38.5}}, {{36.3, 37.7}, {36.3, 37.7}}, {{36.4, 38.1}, {38.1}, {38.0}, {36.4, 38.0}}, {{37.2, 38.0}, {37.9}, {37.9}, {37.2, 37.8}}, {{37.0, 37.8}, {37.9}, {37.9}, {37.0, 38.0}}, {{37.6, 38.4}, {38.4}, {37.6, 38.6}}, {{36.5, 38.3}, {36.5, 38.3}}, {{36.8, 38.8}, {38.8}, {38.7}, {38.7}, {36.8, 38.5}}, {{30.0, 36.1}, {30.0, 36.1}}, {{35.9, 38.7, 38.8}, {38.5}, {35.9, 38.5}}, {{21.9, 31.8}, {21.9, 31.8}}, {{41.8, 44.9}, {44.9}, {44.7}, {44.7}, {41.8, 44.5}}, {{42.3, 44.8}, {45.0, 45.3, 45.5}, {45.1, 45.2}, {44.9}, {45.0}, {45.0}, {44.9}, {45.0, 45.2}, {42.3, 45.3, 45.6}};
		}
	}
}
