netcdf mask {
	:date_created = "20200811T114628";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200811T114628";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 13;
			channels = 4;
			categories = 52;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  81.1, 60.6, 65.7, 75.6, 68.9, 76.1, 75.9, 46.7, 71.2, 76.3, 76.3, 91.4, 60.0;
			max_depth =  87.6, 65.4, 69.2, 78.4, 74.4, 80.2, 81.1, 51.6, 74.9, 91.3, 91.2, 93.9, 63.6;
			start_time = 129179012638710144, 129179010193241472, 129179008324491392, 129179010969022720, 129179014284022656, 129179013662460160, 129179014450585088, 129179012297460224, 129179015636835200, 129179019049335168, 129179019207772672, 129179019252460160, 129179007918085120;
			end_time = 129179012687460096, 129179010278397696, 129179008352772736, 129179010997460096, 129179014328710144, 129179013699022592, 129179014483085184, 129179012325897600, 129179015661210112, 129179019130585216, 129179019264647680, 129179019431210112, 129179007954647680;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "27", "27", "27", "27", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "0", "0", "0", "0", "27", "27", "27", "27";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "120", "200";
			region_channels = 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15;
			mask_times = {1.291790126387101e+17, 1.291790126427727e+17, 1.291790126468351e+17, 1.291790126508977e+17, 1.291790126549603e+17, 1.291790126590226e+17, 1.291790126630852e+17, 1.291790126671476e+17, 1.291790126712101e+17, 1.291790126752727e+17, 1.291790126793352e+17, 1.291790126833976e+17, 1.291790126874601e+17},
			             {1.291790101932415e+17, 1.291790101971476e+17, 1.291790102012102e+17, 1.291790102052726e+17, 1.291790102093352e+17, 1.291790102133978e+17, 1.291790102174601e+17, 1.291790102215227e+17, 1.291790102255852e+17, 1.291790102296476e+17, 1.291790102337102e+17, 1.291790102377727e+17, 1.291790102418351e+17, 1.291790102458976e+17, 1.291790102499602e+17, 1.291790102540227e+17, 1.291790102580851e+17, 1.291790102621476e+17, 1.291790102662102e+17, 1.291790102702726e+17, 1.291790102743352e+17, 1.291790102783977e+17},
			             {1.291790083244914e+17, 1.291790083283977e+17, 1.291790083324602e+17, 1.291790083365226e+17, 1.291790083405852e+17, 1.291790083446477e+17, 1.291790083487101e+17, 1.291790083527727e+17},
			             {1.291790109690227e+17, 1.291790109729289e+17, 1.291790109769915e+17, 1.291790109812102e+17, 1.291790109852726e+17, 1.291790109893352e+17, 1.291790109933978e+17, 1.291790109974601e+17},
			             {1.291790142840227e+17, 1.291790142880851e+17, 1.291790142921477e+17, 1.291790142962102e+17, 1.291790143002726e+17, 1.291790143043352e+17, 1.291790143083976e+17, 1.291790143124602e+17, 1.291790143165228e+17, 1.291790143205851e+17, 1.291790143246477e+17, 1.291790143287101e+17},
			             {1.291790136624602e+17, 1.291790136665226e+17, 1.291790136705852e+17, 1.291790136746477e+17, 1.291790136787103e+17, 1.291790136827727e+17, 1.291790136868351e+17, 1.291790136908977e+17, 1.291790136949603e+17, 1.291790136990226e+17},
			             {1.291790144505851e+17, 1.291790144546477e+17, 1.291790144587103e+17, 1.291790144627726e+17, 1.291790144668352e+17, 1.291790144708977e+17, 1.291790144749603e+17, 1.291790144790227e+17, 1.291790144830852e+17},
			             {1.291790122974602e+17, 1.291790123015227e+17, 1.291790123055852e+17, 1.291790123096476e+17, 1.291790123137102e+17, 1.291790123177727e+17, 1.291790123218351e+17, 1.291790123258976e+17},
			             {1.291790156368352e+17, 1.291790156408977e+17, 1.291790156449601e+17, 1.291790156490226e+17, 1.291790156530852e+17, 1.291790156571476e+17, 1.291790156612101e+17},
			             {1.291790190493352e+17, 1.291790190533976e+17, 1.291790190574602e+17, 1.291790190615227e+17, 1.291790190655852e+17, 1.291790190696476e+17, 1.291790190737101e+17, 1.291790190777727e+17, 1.291790190818353e+17, 1.291790190858977e+17, 1.291790190899602e+17, 1.291790190940227e+17, 1.291790190980852e+17, 1.291790191021476e+17, 1.291790191062102e+17, 1.291790191102728e+17, 1.291790191143351e+17, 1.291790191183977e+17, 1.291790191224603e+17, 1.291790191265226e+17, 1.291790191305852e+17},
			             {1.291790192077727e+17, 1.291790192118351e+17, 1.291790192158977e+17, 1.291790192199602e+17, 1.291790192240227e+17, 1.291790192280852e+17, 1.291790192319914e+17, 1.291790192362102e+17, 1.291790192402728e+17, 1.291790192443351e+17, 1.291790192483977e+17, 1.291790192524602e+17, 1.291790192565226e+17, 1.291790192605852e+17, 1.291790192646477e+17},
			             {1.291790192524602e+17, 1.291790192565226e+17, 1.291790192605852e+17, 1.291790192646477e+17, 1.291790192687101e+17, 1.291790192727726e+17, 1.291790192768352e+17, 1.291790192808977e+17, 1.291790192849601e+17, 1.291790192890227e+17, 1.291790192930852e+17, 1.291790192971476e+17, 1.291790193012102e+17, 1.291790193052727e+17, 1.291790193091789e+17, 1.291790193133976e+17, 1.291790193174602e+17, 1.291790193215227e+17, 1.291790193255852e+17, 1.291790193296476e+17, 1.291790193337101e+17, 1.291790193377727e+17, 1.291790193418353e+17, 1.291790193458976e+17, 1.291790193499602e+17, 1.291790193540227e+17, 1.291790193580852e+17, 1.291790193621476e+17, 1.291790193662102e+17, 1.291790193702728e+17, 1.291790193743351e+17, 1.291790193783977e+17, 1.291790193824603e+17, 1.291790193865226e+17, 1.291790193905852e+17, 1.291790193944914e+17, 1.291790193987101e+17, 1.291790194027727e+17, 1.291790194068352e+17, 1.291790194108977e+17, 1.291790194149601e+17, 1.291790194190227e+17, 1.291790194229289e+17, 1.291790194271476e+17, 1.291790194312101e+17},
			             {1.291790079180851e+17, 1.291790079221476e+17, 1.291790079262102e+17, 1.291790079302726e+17, 1.291790079343351e+17, 1.291790079383977e+17, 1.291790079424602e+17, 1.291790079465226e+17, 1.291790079505852e+17, 1.291790079546477e+17};
			mask_depths = {{81.1, 87.6}, {81.1, 87.6}, {81.1, 87.6}, {81.1, 87.6}, {81.1, 87.6}, {81.1, 87.6}, {81.1, 87.6}, {81.1, 87.5}, {81.1, 87.5}, {81.1, 87.5}, {81.1, 87.5}, {81.1, 87.5}, {81.1, 87.4}}, {{60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}, {60.6, 65.4}}, {{65.7, 69.2}, {65.7, 69.2}, {65.7, 69.2}, {65.7, 69.2}, {65.7, 69.2}, {65.7, 69.2}, {65.7, 69.2}, {65.7, 69.2}}, {{75.6, 78.4}, {75.6, 78.4}, {75.6, 78.4}, {75.6, 78.4}, {75.6, 78.4}, {75.6, 78.4}, {75.6, 78.4}, {75.6, 78.4}}, {{68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}, {68.9, 74.4}}, {{76.1, 80.2}, {76.1, 80.2}, {76.1, 80.2}, {76.1, 80.2}, {76.1, 80.2}, {76.1, 80.2}, {76.1, 80.2}, {76.1, 80.2}, {76.1, 80.2}, {76.1, 80.2}}, {{75.9, 81.1}, {75.9, 81.1}, {75.9, 81.1}, {75.9, 81.1}, {75.9, 81.1}, {75.9, 81.1}, {75.9, 81.1}, {75.9, 81.1}, {75.9, 81.1}}, {{46.7, 51.6}, {46.7, 51.6}, {46.7, 51.6}, {46.7, 51.6}, {46.7, 51.6}, {46.7, 51.6}, {46.7, 51.6}, {46.7, 51.6}}, {{71.2, 74.9}, {71.2, 74.9}, {71.2, 74.9}, {71.2, 74.9}, {71.2, 74.9}, {71.2, 74.9}, {71.2, 74.9}}, {{76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}, {76.3, 91.3}}, {{76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}, {76.3, 91.2}}, {{91.4, 93.1}, {91.4, 93.1}, {91.4, 93.1}, {91.4, 93.1}, {91.4, 93.1}, {91.4, 93.1}, {91.4, 93.1}, {91.4, 93.2}, {91.4, 93.3}, {91.4, 93.3}, {91.4, 93.3}, {91.4, 93.3}, {91.4, 93.3}, {91.4, 93.4}, {91.4, 93.4}, {91.4, 93.4}, {91.4, 93.5}, {91.4, 93.5}, {91.4, 93.5}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.6}, {91.4, 93.7}, {91.4, 93.7}, {91.4, 93.8}, {91.4, 93.8}, {91.4, 93.8}, {91.4, 93.8}, {91.4, 93.9}, {91.4, 93.9}, {91.4, 93.9}, {91.4, 93.9}, {91.4, 93.9}, {91.4, 93.9}, {91.4, 93.9}, {91.4, 93.9}}, {{60.0, 60.0, 63.6, 63.6}, {60.0, 63.6}, {60.0, 63.6}, {60.0, 63.6}, {60.0, 63.6}, {60.0, 63.6}, {60.0, 63.6}, {60.0, 63.6}, {60.0, 63.6}, {60.0, 63.6}};
		}
	}
}
