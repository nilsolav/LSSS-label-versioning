netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 2;
			channels = 4;
			categories = 8;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0, 46.8;
			max_depth =  57.0, 54.6;
			start_time = 129162930133164032, 129162944163945344;
			end_time = 129162955602382848, 129162944276601600;
			region_id = 1, 2;
			region_name = "Layer1","Layer1";
			region_provenance = "LSSS", "LSSS";
			region_comment = "", "";
			region_category_names = "0", "0", "0", "0", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1, 2, 3, 4, 5, 6, 7, 8;
			region_type = analysis, analysis;
			channel_names = "18", "38", "120", "200";
			region_channels = 15, 15;
			mask_times = {1.29162930133164e+17, 1.29162930136289e+17, 1.291629301395704e+17, 1.291629301426953e+17, 1.291629301459766e+17, 1.291629301492579e+17, 1.291629301523828e+17, 1.29162930155664e+17, 1.291629301587891e+17, 1.291629301620704e+17, 1.291629301653516e+17, 1.291629301684765e+17, 1.291629301717578e+17, 1.291629301748828e+17, 1.291629301781641e+17, 1.291629301814454e+17, 1.291629301845704e+17, 1.291629301878515e+17, 1.291629301909766e+17, 1.291629301942579e+17, 1.291629301975391e+17, 1.291629302006641e+17, 1.291629302039453e+17, 1.291629302072266e+17, 1.291629302103515e+17, 1.291629302136329e+17, 1.291629302167579e+17, 1.29162930220039e+17, 1.29162930223164e+17, 1.291629302264454e+17, 1.291629302297266e+17, 1.291629302328516e+17, 1.291629302361329e+17, 1.291629302394141e+17, 1.29162930242539e+17, 1.291629302458204e+17, 1.291629302489454e+17, 1.291629302522266e+17, 1.291629302555078e+17, 1.291629302586328e+17, 1.291629302619141e+17, 1.291629302650391e+17, 1.291629302683204e+17, 1.291629302716015e+17, 1.291629302747265e+17, 1.291629302780078e+17, 1.291629302811329e+17, 1.291629302844141e+17, 1.291629302876954e+17, 1.291629302908204e+17, 1.291629302941016e+17, 1.291629302973829e+17, 1.291629303005079e+17, 1.291629303037891e+17, 1.29162930306914e+17, 1.291629303101953e+17, 1.291629303134766e+17, 1.291629303166016e+17, 1.291629303198829e+17, 1.29162930323164e+17, 1.291629303262892e+17, 1.291629303295704e+17, 1.291629303326954e+17, 1.291629303359766e+17, 1.291629303392579e+17, 1.291629303423828e+17, 1.291629303456641e+17, 1.291629303487891e+17, 1.291629303520704e+17, 1.291629303553516e+17, 1.291629303584765e+17, 1.29162930361758e+17, 1.291629303648828e+17, 1.291629303681641e+17, 1.291629303714454e+17, 1.291629303745704e+17, 1.291629303778515e+17, 1.291629303811328e+17, 1.291629303842579e+17, 1.291629303875391e+17, 1.291629303908204e+17, 1.291629303939453e+17, 1.291629303972266e+17, 1.291629304003516e+17, 1.291629304036329e+17, 1.291629304069142e+17, 1.29162930410039e+17, 1.291629304133203e+17, 1.291629304164454e+17, 1.291629304197266e+17, 1.291629304230079e+17, 1.291629304261329e+17, 1.291629304294141e+17, 1.29162930432539e+17, 1.291629304358204e+17, 1.291629304391016e+17, 1.291629304422266e+17, 1.291629304455078e+17, 1.291629304486328e+17, 1.291629304519141e+17, 1.291629304551953e+17, 1.291629304583204e+17, 1.291629304616017e+17, 1.291629304648828e+17, 1.291629304680078e+17, 1.291629304712891e+17, 1.291629304744141e+17, 1.291629304776954e+17, 1.291629304809766e+17, 1.291629304841016e+17, 1.291629304873828e+17, 1.291629304905079e+17, 1.291629304937892e+17, 1.291629304970703e+17, 1.291629305001953e+17, 1.291629305034766e+17, 1.291629305066016e+17, 1.291629305098828e+17, 1.291629305131642e+17, 1.291629305162892e+17, 1.291629305195703e+17, 1.291629305228516e+17, 1.291629305259766e+17, 1.291629305292579e+17, 1.291629305323828e+17, 1.291629305356641e+17, 1.291629305389453e+17, 1.291629305420703e+17, 1.291629305453516e+17, 1.291629305486328e+17, 1.291629305517578e+17, 1.291629305550391e+17, 1.291629305581641e+17, 1.291629305614454e+17, 1.291629305645704e+17, 1.291629305678516e+17, 1.291629305711328e+17, 1.291629305742578e+17, 1.291629305775391e+17, 1.291629305806641e+17, 1.291629305839453e+17, 1.291629305872266e+17, 1.291629305903516e+17, 1.291629305936328e+17, 1.291629305967578e+17, 1.291629306000392e+17, 1.291629306033203e+17, 1.291629306064453e+17, 1.291629306097266e+17, 1.291629306128516e+17, 1.291629306161329e+17, 1.291629306194141e+17, 1.291629306225391e+17, 1.291629306258203e+17, 1.291629306289453e+17, 1.291629306322266e+17, 1.291629306355078e+17, 1.291629306386328e+17, 1.291629306419141e+17, 1.291629306451953e+17, 1.291629306483204e+17, 1.291629306516017e+17, 1.291629306547267e+17, 1.291629306580078e+17, 1.291629306611328e+17, 1.291629306644141e+17, 1.291629306676954e+17, 1.291629306708204e+17, 1.291629306741016e+17, 1.291629306773828e+17, 1.291629306805078e+17, 1.291629306837892e+17, 1.291629306870703e+17, 1.291629306901953e+17, 1.291629306934766e+17, 1.291629306966016e+17, 1.291629306998828e+17, 1.291629307031642e+17, 1.291629307062892e+17, 1.291629307095703e+17, 1.291629307126953e+17, 1.291629307159767e+17, 1.291629307192579e+17, 1.291629307223828e+17, 1.291629307256641e+17, 1.291629307289454e+17, 1.291629307320703e+17, 1.291629307353517e+17, 1.291629307384767e+17, 1.291629307417578e+17, 1.291629307450391e+17, 1.291629307481642e+17, 1.291629307514454e+17, 1.291629307545704e+17, 1.291629307578516e+17, 1.291629307611329e+17, 1.291629307642578e+17, 1.291629307675391e+17, 1.291629307706642e+17, 1.291629307739453e+17, 1.291629307772266e+17, 1.291629307803516e+17, 1.291629307836329e+17, 1.291629307867578e+17, 1.291629307900392e+17, 1.291629307933203e+17, 1.291629307964453e+17, 1.291629307997266e+17, 1.291629308028517e+17, 1.291629308061329e+17, 1.291629308094141e+17, 1.291629308125391e+17, 1.291629308158204e+17, 1.291629308189453e+17, 1.291629308222267e+17, 1.291629308255078e+17, 1.291629308286328e+17, 1.291629308319141e+17, 1.291629308350391e+17, 1.291629308383204e+17, 1.291629308416015e+17, 1.291629308447267e+17, 1.291629308480078e+17, 1.291629308511328e+17, 1.291629308544141e+17, 1.291629308576954e+17, 1.291629308608204e+17, 1.291629308641016e+17, 1.291629308672266e+17, 1.291629308705079e+17, 1.291629308737891e+17, 1.291629308769142e+17, 1.291629308801953e+17, 1.291629308833203e+17, 1.291629308866016e+17, 1.291629308898829e+17, 1.291629308930079e+17, 1.29162930896289e+17, 1.291629308994141e+17, 1.291629309026954e+17, 1.291629309059766e+17, 1.291629309091016e+17, 1.291629309123828e+17, 1.291629309155078e+17, 1.291629309187891e+17, 1.291629309220704e+17, 1.291629309251954e+17, 1.291629309284765e+17, 1.291629309316017e+17, 1.291629309348828e+17, 1.291629309381641e+17, 1.291629309412891e+17, 1.291629309445704e+17, 1.291629309476954e+17, 1.291629309509766e+17, 1.291629309542578e+17, 1.291629309573829e+17, 1.291629309606641e+17, 1.291629309639453e+17, 1.291629309670703e+17, 1.291629309703516e+17, 1.291629309734766e+17, 1.291629309767579e+17, 1.291629309798829e+17, 1.29162930983164e+17, 1.291629309864453e+17, 1.291629309895703e+17, 1.291629309928516e+17, 1.291629309959766e+17, 1.291629309992579e+17, 1.29162931002539e+17, 1.291629310056641e+17, 1.291629310089454e+17, 1.291629310122266e+17, 1.291629310153516e+17, 1.291629310186328e+17, 1.291629310217578e+17, 1.291629310250391e+17, 1.291629310283204e+17, 1.291629310314454e+17, 1.291629310347265e+17, 1.291629310378516e+17, 1.291629310411328e+17, 1.291629310444141e+17, 1.291629310475391e+17, 1.291629310508204e+17, 1.291629310539453e+17, 1.291629310572266e+17, 1.291629310605079e+17, 1.291629310636329e+17, 1.29162931066914e+17, 1.291629310701955e+17, 1.291629310733203e+17, 1.291629310766016e+17, 1.291629310797266e+17, 1.291629310830079e+17, 1.291629310861329e+17, 1.29162931089414e+17, 1.291629310926954e+17, 1.291629310958203e+17, 1.291629310991016e+17, 1.291629311023828e+17, 1.291629311055078e+17, 1.29162931108789e+17, 1.291629311119141e+17, 1.291629311151954e+17, 1.291629311183204e+17, 1.291629311216015e+17, 1.291629311248829e+17, 1.291629311280078e+17, 1.291629311312891e+17, 1.291629311344141e+17, 1.291629311376954e+17, 1.291629311409765e+17, 1.291629311441015e+17, 1.291629311473829e+17, 1.291629311506641e+17, 1.291629311537891e+17, 1.291629311570705e+17, 1.291629311601953e+17, 1.291629311634766e+17, 1.291629311666016e+17, 1.291629311698829e+17, 1.29162931173164e+17, 1.29162931176289e+17, 1.291629311795704e+17, 1.291629311826953e+17, 1.291629311859766e+17, 1.291629311892579e+17, 1.291629311923828e+17, 1.29162931195664e+17, 1.291629311989454e+17, 1.291629312020704e+17, 1.291629312053516e+17, 1.291629312084765e+17, 1.29162931211758e+17, 1.291629312148828e+17, 1.291629312181641e+17, 1.291629312214454e+17, 1.291629312245704e+17, 1.291629312278515e+17, 1.291629312309765e+17, 1.291629312342579e+17, 1.291629312375391e+17, 1.291629312406641e+17, 1.291629312439453e+17, 1.291629312472266e+17, 1.291629312503515e+17, 1.291629312536329e+17, 1.291629312567579e+17, 1.29162931260039e+17, 1.29162931263164e+17, 1.291629312664454e+17, 1.291629312697266e+17, 1.291629312728516e+17, 1.291629312761329e+17, 1.291629312792579e+17, 1.29162931282539e+17, 1.291629312858204e+17, 1.291629312889454e+17, 1.291629312922266e+17, 1.291629312955078e+17, 1.29162931298633e+17, 1.291629313019141e+17, 1.291629313050391e+17, 1.291629313083204e+17, 1.291629313116017e+17, 1.291629313147265e+17, 1.291629313180079e+17, 1.291629313211329e+17, 1.291629313244141e+17, 1.291629313276954e+17, 1.291629313308204e+17, 1.291629313341016e+17, 1.291629313372265e+17, 1.291629313405079e+17, 1.291629313436329e+17, 1.29162931346914e+17, 1.291629313501953e+17, 1.291629313533204e+17, 1.291629313566016e+17, 1.291629313598829e+17, 1.291629313630079e+17, 1.291629313662892e+17, 1.291629313695703e+17, 1.291629313726954e+17, 1.291629313759766e+17, 1.291629313791016e+17, 1.291629313823828e+17, 1.291629313855078e+17, 1.291629313887891e+17, 1.291629313920704e+17, 1.291629313951954e+17, 1.291629313984765e+17, 1.291629314016015e+17, 1.291629314048828e+17, 1.291629314081641e+17, 1.291629314112891e+17, 1.291629314145704e+17, 1.291629314176954e+17, 1.291629314209766e+17, 1.291629314242579e+17, 1.291629314273829e+17, 1.291629314306641e+17, 1.291629314337891e+17, 1.291629314370703e+17, 1.291629314403516e+17, 1.291629314434766e+17, 1.291629314467579e+17, 1.29162931450039e+17, 1.291629314531642e+17, 1.291629314564453e+17, 1.291629314595704e+17, 1.291629314628516e+17, 1.291629314661329e+17, 1.291629314692579e+17, 1.291629314725391e+17, 1.291629314756641e+17, 1.291629314789454e+17, 1.291629314822266e+17, 1.291629314853516e+17, 1.291629314886328e+17, 1.291629314919141e+17, 1.291629314950391e+17, 1.291629314983204e+17, 1.291629315014454e+17, 1.291629315047265e+17, 1.291629315080078e+17, 1.291629315111329e+17, 1.291629315144141e+17, 1.291629315175391e+17, 1.291629315208204e+17, 1.291629315241016e+17, 1.291629315272266e+17, 1.291629315305078e+17, 1.291629315336329e+17, 1.29162931536914e+17, 1.291629315401953e+17, 1.291629315433203e+17, 1.291629315466016e+17, 1.291629315497266e+17, 1.291629315530079e+17, 1.291629315562892e+17, 1.291629315594141e+17, 1.291629315626953e+17, 1.291629315658204e+17, 1.291629315691016e+17, 1.291629315723828e+17, 1.291629315755078e+17, 1.291629315787891e+17, 1.291629315819141e+17, 1.291629315851954e+17, 1.291629315884767e+17, 1.291629315916015e+17, 1.291629315948828e+17, 1.291629315980079e+17, 1.291629316012891e+17, 1.291629316045702e+17, 1.291629316076954e+17, 1.291629316109766e+17, 1.291629316141016e+17, 1.291629316173828e+17, 1.291629316205079e+17, 1.291629316237891e+17, 1.291629316270703e+17, 1.291629316301953e+17, 1.291629316334766e+17, 1.291629316366016e+17, 1.291629316398829e+17, 1.291629316431642e+17, 1.29162931646289e+17, 1.291629316495703e+17, 1.291629316528516e+17, 1.291629316559766e+17, 1.291629316592577e+17, 1.291629316623828e+17, 1.291629316656641e+17, 1.291629316689453e+17, 1.291629316720703e+17, 1.291629316753517e+17, 1.291629316784765e+17, 1.291629316817578e+17, 1.291629316850391e+17, 1.291629316881641e+17, 1.291629316914452e+17, 1.291629316945704e+17, 1.291629316978516e+17, 1.291629317011328e+17, 1.291629317042578e+17, 1.291629317075391e+17, 1.291629317106641e+17, 1.291629317139453e+17, 1.291629317172266e+17, 1.291629317203516e+17, 1.291629317236328e+17, 1.291629317267579e+17, 1.291629317300392e+17, 1.291629317333203e+17, 1.291629317364453e+17, 1.291629317397266e+17, 1.291629317430079e+17, 1.291629317461327e+17, 1.291629317494141e+17, 1.291629317525391e+17, 1.291629317558203e+17, 1.291629317591016e+17, 1.291629317622267e+17, 1.291629317655078e+17, 1.291629317686328e+17, 1.291629317719141e+17, 1.291629317751954e+17, 1.291629317783203e+17, 1.291629317816017e+17, 1.291629317847267e+17, 1.291629317880078e+17, 1.291629317912891e+17, 1.291629317944141e+17, 1.291629317976954e+17, 1.291629318008204e+17, 1.291629318041016e+17, 1.291629318073828e+17, 1.291629318105078e+17, 1.291629318137891e+17, 1.291629318169142e+17, 1.291629318201953e+17, 1.291629318234766e+17, 1.291629318266016e+17, 1.291629318298829e+17, 1.291629318330077e+17, 1.291629318362892e+17, 1.291629318395703e+17, 1.291629318426953e+17, 1.291629318459766e+17, 1.291629318491017e+17, 1.291629318523828e+17, 1.291629318556641e+17, 1.291629318587891e+17, 1.291629318620704e+17, 1.291629318651953e+17, 1.291629318684767e+17, 1.291629318717578e+17, 1.291629318748828e+17, 1.291629318781641e+17, 1.291629318812891e+17, 1.291629318845704e+17, 1.291629318878516e+17, 1.291629318909766e+17, 1.291629318942578e+17, 1.291629318973828e+17, 1.291629319006641e+17, 1.291629319039453e+17, 1.291629319070703e+17, 1.291629319103516e+17, 1.291629319134766e+17, 1.291629319167579e+17, 1.291629319200392e+17, 1.291629319231642e+17, 1.291629319264453e+17, 1.291629319295703e+17, 1.291629319328516e+17, 1.291629319361329e+17, 1.291629319392579e+17, 1.291629319425391e+17, 1.291629319456641e+17, 1.291629319489453e+17, 1.291629319522267e+17, 1.291629319553516e+17, 1.291629319586328e+17, 1.291629319617578e+17, 1.291629319650391e+17, 1.291629319683204e+17, 1.291629319714454e+17, 1.291629319747267e+17, 1.291629319778516e+17, 1.291629319811328e+17, 1.291629319844142e+17, 1.291629319875391e+17, 1.291629319908204e+17, 1.291629319941016e+17, 1.291629319972266e+17, 1.291629320005078e+17, 1.291629320036329e+17, 1.291629320069142e+17, 1.291629320101953e+17, 1.291629320133203e+17, 1.291629320166016e+17, 1.291629320198829e+17, 1.291629320230079e+17, 1.291629320262892e+17, 1.291629320294141e+17, 1.291629320326953e+17, 1.291629320359766e+17, 1.291629320391017e+17, 1.291629320423828e+17, 1.291629320456641e+17, 1.291629320487891e+17, 1.291629320520704e+17, 1.291629320551953e+17, 1.291629320584767e+17, 1.291629320616017e+17, 1.291629320648828e+17, 1.291629320681641e+17, 1.291629320712891e+17, 1.291629320745704e+17, 1.291629320776954e+17, 1.291629320809766e+17, 1.291629320842579e+17, 1.291629320873828e+17, 1.291629320906641e+17, 1.291629320939453e+17, 1.291629320970703e+17, 1.291629321003516e+17, 1.291629321034766e+17, 1.291629321067579e+17, 1.29162932110039e+17, 1.291629321131642e+17, 1.291629321164453e+17, 1.291629321195703e+17, 1.291629321228516e+17, 1.291629321261329e+17, 1.291629321292579e+17, 1.29162932132539e+17, 1.291629321356641e+17, 1.291629321389454e+17, 1.291629321422266e+17, 1.291629321453516e+17, 1.291629321486328e+17, 1.291629321517578e+17, 1.291629321550391e+17, 1.291629321583204e+17, 1.291629321614454e+17, 1.291629321647265e+17, 1.291629321680078e+17, 1.291629321711329e+17, 1.291629321744141e+17, 1.291629321775391e+17, 1.291629321808204e+17, 1.291629321841016e+17, 1.291629321872266e+17, 1.291629321905079e+17, 1.291629321936329e+17, 1.29162932196914e+17, 1.291629322001953e+17, 1.291629322033203e+17, 1.291629322066016e+17, 1.291629322097266e+17, 1.291629322130079e+17, 1.291629322161329e+17, 1.29162932219414e+17, 1.291629322226953e+17, 1.291629322258204e+17, 1.291629322291016e+17, 1.291629322323828e+17, 1.291629322355078e+17, 1.291629322387891e+17, 1.291629322419141e+17, 1.291629322451954e+17, 1.291629322483204e+17, 1.291629322516015e+17, 1.291629322548828e+17, 1.291629322580078e+17, 1.291629322612891e+17, 1.291629322644141e+17, 1.291629322676954e+17, 1.291629322709766e+17, 1.291629322741016e+17, 1.291629322773829e+17, 1.291629322805079e+17, 1.291629322837891e+17, 1.291629322870703e+17, 1.291629322901953e+17, 1.291629322934766e+17, 1.291629322966016e+17, 1.291629322998829e+17, 1.29162932303164e+17, 1.29162932306289e+17, 1.291629323095703e+17, 1.291629323126954e+17, 1.291629323159766e+17, 1.291629323192579e+17, 1.291629323223828e+17, 1.291629323256641e+17, 1.291629323287891e+17, 1.291629323320704e+17, 1.291629323353516e+17, 1.291629323384765e+17, 1.291629323417578e+17, 1.291629323448828e+17, 1.291629323481641e+17, 1.291629323514454e+17, 1.291629323545704e+17, 1.291629323578515e+17, 1.291629323611329e+17, 1.291629323642578e+17, 1.291629323675391e+17, 1.291629323706641e+17, 1.291629323739453e+17, 1.291629323772265e+17, 1.291629323803516e+17, 1.291629323836329e+17, 1.29162932386914e+17, 1.29162932390039e+17, 1.291629323933204e+17, 1.291629323964453e+17, 1.291629323997266e+17, 1.291629324030079e+17, 1.291629324061329e+17, 1.29162932409414e+17, 1.291629324125391e+17, 1.291629324158204e+17, 1.291629324189454e+17, 1.291629324222266e+17, 1.29162932425508e+17, 1.291629324286328e+17, 1.291629324319141e+17, 1.291629324351954e+17, 1.291629324383204e+17, 1.291629324416015e+17, 1.291629324447265e+17, 1.291629324480079e+17, 1.291629324511328e+17, 1.291629324544141e+17, 1.291629324576954e+17, 1.291629324608204e+17, 1.291629324641015e+17, 1.291629324673829e+17, 1.291629324705079e+17, 1.291629324737891e+17, 1.29162932476914e+17, 1.291629324801955e+17, 1.291629324834766e+17, 1.291629324866016e+17, 1.291629324898829e+17, 1.291629324930079e+17, 1.29162932496289e+17, 1.291629324995704e+17, 1.291629325026954e+17, 1.291629325059766e+17, 1.291629325091016e+17, 1.291629325123828e+17, 1.291629325156641e+17, 1.29162932518789e+17, 1.291629325220704e+17, 1.291629325251954e+17, 1.291629325284765e+17, 1.291629325317578e+17, 1.291629325348829e+17, 1.291629325381641e+17, 1.291629325412891e+17, 1.291629325445704e+17, 1.291629325478516e+17, 1.291629325509765e+17, 1.291629325542579e+17, 1.291629325573829e+17, 1.291629325606641e+17, 1.291629325639453e+17, 1.291629325670705e+17, 1.291629325703516e+17, 1.291629325734766e+17, 1.291629325767579e+17, 1.291629325800392e+17, 1.29162932583164e+17, 1.291629325864454e+17, 1.291629325895704e+17, 1.291629325928516e+17, 1.291629325961329e+17, 1.291629325992579e+17, 1.291629326025391e+17, 1.29162932605664e+17, 1.291629326089454e+17, 1.291629326122266e+17, 1.291629326153516e+17, 1.291629326186328e+17, 1.29162932621758e+17, 1.291629326250391e+17, 1.291629326283204e+17, 1.291629326314454e+17, 1.291629326347267e+17, 1.291629326378515e+17, 1.291629326411329e+17, 1.291629326442579e+17, 1.291629326475391e+17, 1.291629326508204e+17, 1.291629326539453e+17, 1.291629326572266e+17, 1.291629326605079e+17, 1.291629326636329e+17, 1.29162932666914e+17, 1.29162932670039e+17, 1.291629326733204e+17, 1.291629326766016e+17, 1.291629326797266e+17, 1.291629326830079e+17, 1.291629326861329e+17, 1.291629326894141e+17, 1.291629326926953e+17, 1.291629326958204e+17, 1.291629326991016e+17, 1.291629327023828e+17, 1.291629327055078e+17, 1.291629327087891e+17, 1.291629327119141e+17, 1.291629327151954e+17, 1.291629327184765e+17, 1.291629327216017e+17, 1.291629327248828e+17, 1.291629327280079e+17, 1.291629327312891e+17, 1.291629327345704e+17, 1.291629327376954e+17, 1.291629327409766e+17, 1.291629327442578e+17, 1.291629327473829e+17, 1.291629327506641e+17, 1.291629327537891e+17, 1.291629327570703e+17, 1.291629327601953e+17, 1.291629327634766e+17, 1.291629327667578e+17, 1.291629327698829e+17, 1.29162932773164e+17, 1.291629327764453e+17, 1.291629327795703e+17, 1.291629327828516e+17, 1.291629327859766e+17, 1.291629327892579e+17, 1.291629327923828e+17, 1.291629327956641e+17, 1.291629327989453e+17, 1.291629328020704e+17, 1.291629328053516e+17, 1.291629328086328e+17, 1.291629328117578e+17, 1.291629328150391e+17, 1.291629328181641e+17, 1.291629328214454e+17, 1.291629328245704e+17, 1.291629328278516e+17, 1.291629328311328e+17, 1.291629328342579e+17, 1.291629328375391e+17, 1.291629328406641e+17, 1.291629328439453e+17, 1.291629328472266e+17, 1.291629328503516e+17, 1.291629328536328e+17, 1.291629328567579e+17, 1.29162932860039e+17, 1.291629328633203e+17, 1.291629328664453e+17, 1.291629328697266e+17, 1.291629328728516e+17, 1.291629328761329e+17, 1.291629328794141e+17, 1.291629328825391e+17, 1.291629328858203e+17, 1.291629328889454e+17, 1.291629328922266e+17, 1.291629328955078e+17, 1.291629328986328e+17, 1.291629329019141e+17, 1.291629329050391e+17, 1.291629329083203e+17, 1.291629329116017e+17, 1.291629329147265e+17, 1.291629329180078e+17, 1.291629329211328e+17, 1.291629329244141e+17, 1.291629329276952e+17, 1.291629329308204e+17, 1.291629329341016e+17, 1.291629329372266e+17, 1.291629329405078e+17, 1.291629329437892e+17, 1.29162932946914e+17, 1.291629329501953e+17, 1.291629329533203e+17, 1.291629329566016e+17, 1.291629329598828e+17, 1.291629329630079e+17, 1.291629329662892e+17, 1.291629329694141e+17, 1.291629329726953e+17, 1.291629329759767e+17, 1.291629329791016e+17, 1.291629329823828e+17, 1.291629329855078e+17, 1.291629329887891e+17, 1.291629329920703e+17, 1.291629329951953e+17, 1.291629329984767e+17, 1.291629330016015e+17, 1.291629330048828e+17, 1.291629330081641e+17, 1.291629330112891e+17, 1.291629330145702e+17, 1.291629330176954e+17, 1.291629330209766e+17, 1.291629330242578e+17, 1.291629330273828e+17, 1.291629330306642e+17, 1.291629330337891e+17, 1.291629330370703e+17, 1.291629330403516e+17, 1.291629330434766e+17, 1.291629330467578e+17, 1.291629330498829e+17, 1.291629330531642e+17, 1.291629330564453e+17, 1.291629330595703e+17, 1.291629330628516e+17, 1.291629330659766e+17, 1.291629330692577e+17, 1.291629330725391e+17, 1.291629330756641e+17, 1.291629330789453e+17, 1.291629330820703e+17, 1.291629330853517e+17, 1.291629330886328e+17, 1.291629330917578e+17, 1.291629330950391e+17, 1.291629330981641e+17, 1.291629331014452e+17, 1.291629331047267e+17, 1.291629331078516e+17, 1.291629331111328e+17, 1.291629331142578e+17, 1.291629331175392e+17, 1.291629331208204e+17, 1.291629331239453e+17, 1.291629331272266e+17, 1.291629331303516e+17, 1.291629331336328e+17, 1.291629331367579e+17, 1.291629331400392e+17, 1.291629331433203e+17, 1.291629331464453e+17, 1.291629331497266e+17, 1.291629331530079e+17, 1.291629331561327e+17, 1.291629331594141e+17, 1.291629331625391e+17, 1.291629331658203e+17, 1.291629331691016e+17, 1.291629331722267e+17, 1.291629331755078e+17, 1.291629331786328e+17, 1.291629331819141e+17, 1.291629331851954e+17, 1.291629331883203e+17, 1.291629331916017e+17, 1.291629331947267e+17, 1.291629331980078e+17, 1.291629332012891e+17, 1.291629332044141e+17, 1.291629332076954e+17, 1.291629332108204e+17, 1.291629332141016e+17, 1.291629332173828e+17, 1.291629332205078e+17, 1.291629332237892e+17, 1.291629332269142e+17, 1.291629332301953e+17, 1.291629332334766e+17, 1.291629332366016e+17, 1.291629332398829e+17, 1.291629332430077e+17, 1.291629332462892e+17, 1.291629332495703e+17, 1.291629332526953e+17, 1.291629332559766e+17, 1.291629332591017e+17, 1.291629332623828e+17, 1.291629332656641e+17, 1.291629332687891e+17, 1.291629332720704e+17, 1.291629332751953e+17, 1.291629332784767e+17, 1.291629332817578e+17, 1.291629332848828e+17, 1.291629332881641e+17, 1.291629332912891e+17, 1.291629332945704e+17, 1.291629332978516e+17, 1.291629333009766e+17, 1.291629333042578e+17, 1.291629333073828e+17, 1.291629333106641e+17, 1.291629333139453e+17, 1.291629333170703e+17, 1.291629333203516e+17, 1.291629333236328e+17, 1.291629333267579e+17, 1.291629333300392e+17, 1.291629333333203e+17, 1.291629333364453e+17, 1.291629333397266e+17, 1.291629333428516e+17, 1.291629333461329e+17, 1.291629333492579e+17, 1.291629333525391e+17, 1.291629333558203e+17, 1.291629333589453e+17, 1.291629333622267e+17, 1.291629333655078e+17, 1.291629333686328e+17, 1.291629333719141e+17, 1.291629333750391e+17, 1.291629333783204e+17, 1.291629333816015e+17, 1.291629333847267e+17, 1.291629333880078e+17, 1.291629333911328e+17, 1.291629333944141e+17, 1.291629333976954e+17, 1.291629334008204e+17, 1.291629334041016e+17, 1.291629334073829e+17, 1.291629334105078e+17, 1.291629334137891e+17, 1.291629334169142e+17, 1.291629334201953e+17, 1.291629334234766e+17, 1.291629334266016e+17, 1.291629334298829e+17, 1.291629334330079e+17, 1.291629334362892e+17, 1.291629334395704e+17, 1.291629334426953e+17, 1.291629334459766e+17, 1.291629334492579e+17, 1.291629334523828e+17, 1.29162933455664e+17, 1.291629334587891e+17, 1.291629334620704e+17, 1.291629334653516e+17, 1.291629334684765e+17, 1.291629334717578e+17, 1.291629334748828e+17, 1.291629334781641e+17, 1.291629334814454e+17, 1.291629334845704e+17, 1.291629334878515e+17, 1.291629334911328e+17, 1.291629334942579e+17, 1.291629334975391e+17, 1.291629335006641e+17, 1.291629335039453e+17, 1.291629335070703e+17, 1.291629335103516e+17, 1.291629335136329e+17, 1.291629335167579e+17, 1.29162933520039e+17, 1.291629335231642e+17, 1.291629335264454e+17, 1.291629335297266e+17, 1.291629335328516e+17, 1.291629335361329e+17, 1.291629335394141e+17, 1.29162933542539e+17, 1.291629335458204e+17, 1.291629335489454e+17, 1.291629335522266e+17, 1.291629335555078e+17, 1.291629335586328e+17, 1.291629335619141e+17, 1.291629335650391e+17, 1.291629335683204e+17, 1.291629335714454e+17, 1.291629335747265e+17, 1.291629335780078e+17, 1.291629335811329e+17, 1.291629335844141e+17, 1.291629335876954e+17, 1.291629335908204e+17, 1.291629335941016e+17, 1.291629335972266e+17, 1.291629336005079e+17, 1.291629336036329e+17, 1.29162933606914e+17, 1.291629336101953e+17, 1.291629336133203e+17, 1.291629336166016e+17, 1.291629336198829e+17, 1.291629336230079e+17, 1.29162933626289e+17, 1.29162933629414e+17, 1.291629336326954e+17, 1.291629336358204e+17, 1.291629336391016e+17, 1.291629336423828e+17, 1.291629336455078e+17, 1.291629336487891e+17, 1.291629336519141e+17, 1.291629336551954e+17, 1.291629336584765e+17, 1.291629336616015e+17, 1.291629336648828e+17, 1.291629336681641e+17, 1.291629336712891e+17, 1.291629336745704e+17, 1.291629336776954e+17, 1.291629336809766e+17, 1.291629336842579e+17, 1.291629336873829e+17, 1.291629336906641e+17, 1.291629336937891e+17, 1.291629336970703e+17, 1.291629337003516e+17, 1.291629337034766e+17, 1.291629337067579e+17, 1.291629337098829e+17, 1.29162933713164e+17, 1.291629337164454e+17, 1.291629337195703e+17, 1.291629337228516e+17, 1.291629337259766e+17, 1.291629337292579e+17, 1.291629337323828e+17, 1.291629337356641e+17, 1.291629337389454e+17, 1.291629337420704e+17, 1.291629337453516e+17, 1.29162933748633e+17, 1.291629337517578e+17, 1.291629337550391e+17, 1.291629337583204e+17, 1.291629337614454e+17, 1.291629337647265e+17, 1.291629337678515e+17, 1.291629337711329e+17, 1.291629337744141e+17, 1.291629337775391e+17, 1.291629337808204e+17, 1.291629337839453e+17, 1.291629337872266e+17, 1.291629337905079e+17, 1.291629337936329e+17, 1.29162933796914e+17, 1.29162933800039e+17, 1.291629338033204e+17, 1.291629338066016e+17, 1.291629338097266e+17, 1.291629338130079e+17, 1.291629338161329e+17, 1.29162933819414e+17, 1.291629338226954e+17, 1.291629338258204e+17, 1.291629338291016e+17, 1.291629338322266e+17, 1.29162933835508e+17, 1.291629338387891e+17, 1.291629338419141e+17, 1.291629338451954e+17, 1.291629338483204e+17, 1.291629338516015e+17, 1.291629338548828e+17, 1.291629338580079e+17, 1.291629338612891e+17, 1.291629338644141e+17, 1.291629338676954e+17, 1.291629338709766e+17, 1.291629338741015e+17, 1.291629338773829e+17, 1.291629338806641e+17, 1.291629338837891e+17, 1.291629338870703e+17, 1.291629338901955e+17, 1.291629338934766e+17, 1.291629338967579e+17, 1.291629338998829e+17, 1.291629339031642e+17, 1.29162933906289e+17, 1.291629339095704e+17, 1.291629339128516e+17, 1.291629339159766e+17, 1.291629339192579e+17, 1.291629339223828e+17, 1.291629339256641e+17, 1.291629339289453e+17, 1.291629339320704e+17, 1.291629339353517e+17, 1.291629339384765e+17, 1.291629339417578e+17, 1.291629339450391e+17, 1.291629339481641e+17, 1.291629339514454e+17, 1.291629339545704e+17, 1.291629339578516e+17, 1.291629339611328e+17, 1.291629339642579e+17, 1.291629339675391e+17, 1.291629339706641e+17, 1.291629339739453e+17, 1.291629339772266e+17, 1.291629339803516e+17, 1.291629339836329e+17, 1.291629339867579e+17, 1.291629339900392e+17, 1.29162933993164e+17, 1.291629339964454e+17, 1.291629339997266e+17, 1.291629340028516e+17, 1.291629340061329e+17, 1.291629340092579e+17, 1.291629340125391e+17, 1.291629340158203e+17, 1.291629340189454e+17, 1.291629340222266e+17, 1.291629340255078e+17, 1.291629340286328e+17, 1.291629340319141e+17, 1.291629340350391e+17, 1.291629340383204e+17, 1.291629340414454e+17, 1.291629340447267e+17, 1.291629340480078e+17, 1.291629340511329e+17, 1.291629340544141e+17, 1.291629340576954e+17, 1.291629340608204e+17, 1.291629340641016e+17, 1.291629340672266e+17, 1.291629340705078e+17, 1.291629340736329e+17, 1.291629340769142e+17, 1.291629340801953e+17, 1.291629340833203e+17, 1.291629340866016e+17, 1.291629340898829e+17, 1.291629340930079e+17, 1.291629340962892e+17, 1.291629340994141e+17, 1.291629341026953e+17, 1.291629341059766e+17, 1.291629341091016e+17, 1.291629341123828e+17, 1.291629341155078e+17, 1.291629341187891e+17, 1.291629341220703e+17, 1.291629341251954e+17, 1.291629341284765e+17, 1.291629341316017e+17, 1.291629341348828e+17, 1.291629341381641e+17, 1.291629341412891e+17, 1.291629341445704e+17, 1.291629341476954e+17, 1.291629341509766e+17, 1.291629341542578e+17, 1.291629341573828e+17, 1.291629341606641e+17, 1.291629341637891e+17, 1.291629341670703e+17, 1.291629341703516e+17, 1.291629341734766e+17, 1.291629341767578e+17, 1.291629341800392e+17, 1.291629341831642e+17, 1.291629341864453e+17, 1.291629341895703e+17, 1.291629341928516e+17, 1.291629341961329e+17, 1.291629341992579e+17, 1.291629342025391e+17, 1.291629342056641e+17, 1.291629342089453e+17, 1.291629342122267e+17, 1.291629342153516e+17, 1.291629342186328e+17, 1.291629342217578e+17, 1.291629342250391e+17, 1.291629342283203e+17, 1.291629342314454e+17, 1.291629342347267e+17, 1.291629342378516e+17, 1.291629342411328e+17, 1.291629342444142e+17, 1.291629342475391e+17, 1.291629342508204e+17, 1.291629342539453e+17, 1.291629342572266e+17, 1.291629342605078e+17, 1.291629342636328e+17, 1.291629342669142e+17, 1.29162934270039e+17, 1.291629342733203e+17, 1.291629342766016e+17, 1.291629342797266e+17, 1.291629342830077e+17, 1.291629342861329e+17, 1.291629342894141e+17, 1.291629342926953e+17, 1.291629342958203e+17, 1.291629342991017e+17, 1.291629343022266e+17, 1.291629343055078e+17, 1.291629343087891e+17, 1.291629343119141e+17, 1.291629343151953e+17, 1.291629343183203e+17, 1.291629343216017e+17, 1.291629343248828e+17, 1.291629343280078e+17, 1.291629343312891e+17, 1.291629343344141e+17, 1.291629343376954e+17, 1.291629343409766e+17, 1.291629343441016e+17, 1.291629343473828e+17, 1.291629343505078e+17, 1.291629343537892e+17, 1.291629343570703e+17, 1.291629343601953e+17, 1.291629343634766e+17, 1.291629343667579e+17, 1.291629343698828e+17, 1.291629343731642e+17, 1.291629343762892e+17, 1.291629343795703e+17, 1.291629343828516e+17, 1.291629343859767e+17, 1.291629343892579e+17, 1.291629343923828e+17, 1.291629343956641e+17, 1.291629343989454e+17, 1.291629344020703e+17, 1.291629344053517e+17, 1.291629344084767e+17, 1.291629344117578e+17, 1.291629344150391e+17, 1.291629344181641e+17, 1.291629344214454e+17, 1.291629344245702e+17, 1.291629344278516e+17, 1.291629344311328e+17, 1.291629344342578e+17, 1.291629344375391e+17, 1.291629344408204e+17, 1.291629344439453e+17, 1.291629344472266e+17, 1.291629344505078e+17, 1.291629344536329e+17, 1.29162934456914e+17, 1.291629344600392e+17, 1.291629344633203e+17, 1.291629344664453e+17, 1.291629344697266e+17, 1.291629344730079e+17, 1.291629344761329e+17, 1.291629344794141e+17, 1.291629344826953e+17, 1.291629344858204e+17, 1.291629344891016e+17, 1.291629344922267e+17, 1.291629344955078e+17, 1.291629344987891e+17, 1.291629345019141e+17, 1.291629345051954e+17, 1.291629345083204e+17, 1.291629345116017e+17, 1.291629345148828e+17, 1.291629345180078e+17, 1.291629345212891e+17, 1.291629345244141e+17, 1.291629345276954e+17, 1.291629345309765e+17, 1.291629345341016e+17, 1.291629345373828e+17, 1.291629345405079e+17, 1.291629345437891e+17, 1.291629345470703e+17, 1.291629345501953e+17, 1.291629345534766e+17, 1.291629345566016e+17, 1.291629345598829e+17, 1.29162934563164e+17, 1.291629345662892e+17, 1.291629345695703e+17, 1.291629345726953e+17, 1.291629345759766e+17, 1.291629345792579e+17, 1.291629345823828e+17, 1.291629345856641e+17, 1.291629345887891e+17, 1.291629345920703e+17, 1.291629345953516e+17, 1.291629345984767e+17, 1.291629346017578e+17, 1.291629346048828e+17, 1.291629346081641e+17, 1.291629346114454e+17, 1.291629346145704e+17, 1.291629346178515e+17, 1.291629346209766e+17, 1.291629346242578e+17, 1.291629346275391e+17, 1.291629346306641e+17, 1.291629346339453e+17, 1.291629346370703e+17, 1.291629346403516e+17, 1.291629346436329e+17, 1.291629346467579e+17, 1.29162934650039e+17, 1.291629346531642e+17, 1.291629346564453e+17, 1.291629346595703e+17, 1.291629346628516e+17, 1.291629346661329e+17, 1.291629346692579e+17, 1.291629346725391e+17, 1.291629346756641e+17, 1.291629346789453e+17, 1.291629346822266e+17, 1.291629346853517e+17, 1.291629346886328e+17, 1.291629346917578e+17, 1.291629346950391e+17, 1.291629346983204e+17, 1.291629347014454e+17, 1.291629347047265e+17, 1.291629347078516e+17, 1.291629347111328e+17, 1.291629347144141e+17, 1.291629347175391e+17, 1.291629347208204e+17, 1.291629347241015e+17, 1.291629347272266e+17, 1.291629347305079e+17, 1.291629347336328e+17, 1.29162934736914e+17, 1.291629347401953e+17, 1.291629347433203e+17, 1.291629347466016e+17, 1.291629347498829e+17, 1.291629347530079e+17, 1.29162934756289e+17, 1.291629347594141e+17, 1.291629347626954e+17, 1.291629347659766e+17, 1.291629347691016e+17, 1.291629347723828e+17, 1.291629347756641e+17, 1.29162934778789e+17, 1.291629347820704e+17, 1.291629347851954e+17, 1.291629347884765e+17, 1.291629347917578e+17, 1.291629347948829e+17, 1.291629347981641e+17, 1.291629348012891e+17, 1.291629348045704e+17, 1.291629348076954e+17, 1.291629348109765e+17, 1.291629348142579e+17, 1.291629348173829e+17, 1.291629348206641e+17, 1.291629348239453e+17, 1.291629348270703e+17, 1.291629348303516e+17, 1.291629348334765e+17, 1.291629348367579e+17, 1.29162934840039e+17, 1.29162934843164e+17, 1.291629348464453e+17, 1.291629348495704e+17, 1.291629348528516e+17, 1.291629348561329e+17, 1.291629348592579e+17, 1.291629348625391e+17, 1.29162934865664e+17, 1.291629348689454e+17, 1.291629348722266e+17, 1.291629348753516e+17, 1.291629348786328e+17, 1.291629348817578e+17, 1.291629348850391e+17, 1.291629348883204e+17, 1.291629348914454e+17, 1.291629348947265e+17, 1.291629348978515e+17, 1.291629349011329e+17, 1.291629349044141e+17, 1.291629349075391e+17, 1.291629349108204e+17, 1.291629349139453e+17, 1.291629349172266e+17, 1.291629349205079e+17, 1.291629349236329e+17, 1.29162934926914e+17, 1.291629349301953e+17, 1.291629349333203e+17, 1.291629349366016e+17, 1.291629349397266e+17, 1.291629349430079e+17, 1.291629349461329e+17, 1.291629349494141e+17, 1.291629349526954e+17, 1.291629349558204e+17, 1.291629349591016e+17, 1.291629349623828e+17, 1.291629349655078e+17, 1.291629349687891e+17, 1.291629349719141e+17, 1.291629349751954e+17, 1.291629349783204e+17, 1.291629349816015e+17, 1.291629349848829e+17, 1.291629349880078e+17, 1.291629349912891e+17, 1.291629349944141e+17, 1.291629349976954e+17, 1.291629350009765e+17, 1.291629350041016e+17, 1.291629350073829e+17, 1.291629350105079e+17, 1.291629350137891e+17, 1.291629350170703e+17, 1.291629350201953e+17, 1.291629350234766e+17, 1.291629350266016e+17, 1.291629350298829e+17, 1.29162935033164e+17, 1.291629350362892e+17, 1.291629350395704e+17, 1.291629350426954e+17, 1.291629350459766e+17, 1.291629350492579e+17, 1.291629350523828e+17, 1.291629350556641e+17, 1.291629350587891e+17, 1.291629350620704e+17, 1.291629350653516e+17, 1.291629350684765e+17, 1.29162935071758e+17, 1.291629350748828e+17, 1.291629350781641e+17, 1.291629350814454e+17, 1.291629350845704e+17, 1.291629350878515e+17, 1.291629350909766e+17, 1.291629350942579e+17, 1.291629350975391e+17, 1.291629351006641e+17, 1.291629351039453e+17, 1.291629351072266e+17, 1.291629351103516e+17, 1.291629351136329e+17, 1.291629351169142e+17, 1.29162935120039e+17, 1.291629351233203e+17, 1.291629351264454e+17, 1.291629351297266e+17, 1.291629351330079e+17, 1.291629351361329e+17, 1.291629351394141e+17, 1.29162935142539e+17, 1.291629351458204e+17, 1.291629351489454e+17, 1.291629351522266e+17, 1.291629351555078e+17, 1.29162935158633e+17, 1.291629351619141e+17, 1.291629351651953e+17, 1.291629351683204e+17, 1.291629351716017e+17, 1.291629351747265e+17, 1.291629351780078e+17, 1.291629351812891e+17, 1.291629351844141e+17, 1.291629351876954e+17, 1.291629351908204e+17, 1.291629351941016e+17, 1.291629351973828e+17, 1.291629352005079e+17, 1.291629352037892e+17, 1.29162935206914e+17, 1.291629352101953e+17, 1.291629352133204e+17, 1.291629352166016e+17, 1.291629352198829e+17, 1.291629352230079e+17, 1.291629352262892e+17, 1.29162935229414e+17, 1.291629352326953e+17, 1.291629352359766e+17, 1.291629352391016e+17, 1.291629352423828e+17, 1.291629352456641e+17, 1.291629352487891e+17, 1.291629352520703e+17, 1.291629352551954e+17, 1.291629352584767e+17, 1.291629352617578e+17, 1.291629352648828e+17, 1.291629352681641e+17, 1.291629352712891e+17, 1.291629352745704e+17, 1.291629352778516e+17, 1.291629352809766e+17, 1.291629352842578e+17, 1.291629352873829e+17, 1.291629352906641e+17, 1.291629352939453e+17, 1.291629352970703e+17, 1.291629353003516e+17, 1.291629353034766e+17, 1.291629353067578e+17, 1.291629353100392e+17, 1.291629353131642e+17, 1.291629353164453e+17, 1.291629353195703e+17, 1.291629353228516e+17, 1.291629353261329e+17, 1.291629353292579e+17, 1.291629353325391e+17, 1.291629353356641e+17, 1.291629353389453e+17, 1.291629353422266e+17, 1.291629353453517e+17, 1.291629353486328e+17, 1.291629353517578e+17, 1.291629353550391e+17, 1.291629353583204e+17, 1.291629353614454e+17, 1.291629353647267e+17, 1.291629353678516e+17, 1.291629353711328e+17, 1.291629353744141e+17, 1.291629353775391e+17, 1.291629353808204e+17, 1.291629353839453e+17, 1.291629353872266e+17, 1.291629353905078e+17, 1.291629353936328e+17, 1.29162935396914e+17, 1.291629354000392e+17, 1.291629354033203e+17, 1.291629354066016e+17, 1.291629354097266e+17, 1.291629354130079e+17, 1.291629354161329e+17, 1.291629354194141e+17, 1.291629354226953e+17, 1.291629354258203e+17, 1.291629354291016e+17, 1.291629354323828e+17, 1.291629354355078e+17, 1.291629354387891e+17, 1.291629354419141e+17, 1.291629354451953e+17, 1.291629354484767e+17, 1.291629354516017e+17, 1.291629354548828e+17, 1.291629354581642e+17, 1.291629354612891e+17, 1.291629354645704e+17, 1.291629354676954e+17, 1.291629354709766e+17, 1.291629354741016e+17, 1.291629354773828e+17, 1.291629354806642e+17, 1.291629354837891e+17, 1.291629354870703e+17, 1.291629354901953e+17, 1.291629354934766e+17, 1.291629354967578e+17, 1.291629354998829e+17, 1.291629355031642e+17, 1.291629355064453e+17, 1.291629355095703e+17, 1.291629355128517e+17, 1.291629355159766e+17, 1.291629355192579e+17, 1.291629355223828e+17, 1.291629355256641e+17, 1.291629355289453e+17, 1.291629355320703e+17, 1.291629355353517e+17, 1.291629355386328e+17, 1.291629355417578e+17, 1.291629355450391e+17, 1.291629355481641e+17, 1.291629355514452e+17, 1.291629355545704e+17, 1.291629355578516e+17, 1.291629355611328e+17, 1.291629355642578e+17, 1.291629355675392e+17, 1.291629355706641e+17, 1.291629355739453e+17, 1.291629355772266e+17, 1.291629355803516e+17, 1.291629355836328e+17, 1.291629355869142e+17, 1.291629355900392e+17, 1.291629355933203e+17, 1.291629355964453e+17, 1.291629355997267e+17, 1.291629356030079e+17, 1.291629356061329e+17, 1.291629356094141e+17, 1.291629356125391e+17, 1.291629356158203e+17, 1.291629356191017e+17, 1.291629356222267e+17, 1.291629356255078e+17, 1.291629356286328e+17, 1.291629356319141e+17, 1.291629356351954e+17, 1.291629356383203e+17, 1.291629356416017e+17, 1.291629356447267e+17, 1.291629356480078e+17, 1.291629356511328e+17, 1.291629356544142e+17, 1.291629356576954e+17, 1.291629356608204e+17, 1.291629356641016e+17, 1.291629356673829e+17, 1.291629356705078e+17, 1.291629356737892e+17, 1.291629356769142e+17, 1.291629356801953e+17, 1.291629356833203e+17, 1.291629356866016e+17, 1.291629356898829e+17, 1.291629356930077e+17, 1.291629356962892e+17, 1.291629356994141e+17, 1.291629357026953e+17, 1.291629357059766e+17, 1.291629357091017e+17, 1.291629357123828e+17, 1.291629357155078e+17, 1.291629357187891e+17, 1.291629357220704e+17, 1.291629357251953e+17, 1.291629357284767e+17, 1.291629357316017e+17, 1.291629357348828e+17, 1.291629357381641e+17, 1.291629357412892e+17, 1.291629357445704e+17, 1.291629357476954e+17, 1.291629357509766e+17, 1.291629357542579e+17, 1.291629357573828e+17, 1.291629357606642e+17, 1.291629357639453e+17, 1.291629357670703e+17, 1.291629357703516e+17, 1.291629357734766e+17, 1.291629357767579e+17, 1.291629357798828e+17, 1.291629357831642e+17, 1.291629357864453e+17, 1.291629357895703e+17, 1.291629357928516e+17, 1.291629357961329e+17, 1.291629357992579e+17, 1.291629358025391e+17, 1.291629358058203e+17, 1.291629358089454e+17, 1.291629358122266e+17, 1.291629358153517e+17, 1.291629358186328e+17, 1.291629358219141e+17, 1.291629358250391e+17, 1.291629358283204e+17, 1.291629358314454e+17, 1.291629358347267e+17, 1.291629358380078e+17, 1.291629358411328e+17, 1.291629358444141e+17, 1.291629358476954e+17, 1.291629358508204e+17, 1.291629358541015e+17, 1.291629358572266e+17, 1.291629358605079e+17, 1.291629358636329e+17, 1.29162935866914e+17, 1.291629358701953e+17, 1.291629358733203e+17, 1.291629358766016e+17, 1.291629358797266e+17, 1.291629358830079e+17, 1.29162935886289e+17, 1.291629358894141e+17, 1.291629358926953e+17, 1.291629358958204e+17, 1.291629358991016e+17, 1.291629359023828e+17, 1.291629359055078e+17, 1.291629359087891e+17, 1.291629359119141e+17, 1.291629359151954e+17, 1.291629359184765e+17, 1.291629359216017e+17, 1.291629359248828e+17, 1.291629359281641e+17, 1.291629359312891e+17, 1.291629359345704e+17, 1.291629359376954e+17, 1.291629359409765e+17, 1.291629359442579e+17, 1.291629359473828e+17, 1.291629359506641e+17, 1.291629359537891e+17, 1.291629359570703e+17, 1.291629359601953e+17, 1.291629359634766e+17, 1.291629359667579e+17, 1.291629359698829e+17, 1.29162935973164e+17, 1.291629359764454e+17, 1.291629359795703e+17, 1.291629359828516e+17, 1.291629359859766e+17, 1.291629359892579e+17, 1.291629359923828e+17, 1.29162935995664e+17, 1.291629359989454e+17, 1.291629360020704e+17, 1.291629360053516e+17, 1.29162936008633e+17, 1.291629360117578e+17, 1.291629360150391e+17, 1.291629360181641e+17, 1.291629360214454e+17, 1.291629360247265e+17, 1.291629360278515e+17, 1.291629360311329e+17, 1.291629360342578e+17, 1.291629360375391e+17, 1.291629360408204e+17, 1.291629360439453e+17, 1.291629360472265e+17, 1.291629360503516e+17, 1.291629360536329e+17, 1.291629360567579e+17, 1.29162936060039e+17, 1.291629360633204e+17, 1.291629360664453e+17, 1.291629360697266e+17, 1.291629360728516e+17, 1.291629360761329e+17, 1.29162936079414e+17, 1.29162936082539e+17, 1.291629360858204e+17, 1.291629360889453e+17, 1.291629360922266e+17, 1.291629360955078e+17, 1.291629360986328e+17, 1.29162936101914e+17, 1.291629361051954e+17, 1.291629361083204e+17, 1.291629361116015e+17, 1.291629361147265e+17, 1.291629361180079e+17, 1.291629361211328e+17, 1.291629361244141e+17, 1.291629361276954e+17, 1.291629361308204e+17, 1.291629361341015e+17, 1.291629361373829e+17, 1.291629361405079e+17, 1.291629361437891e+17, 1.29162936146914e+17, 1.291629361501955e+17, 1.291629361534766e+17, 1.291629361566016e+17, 1.291629361598829e+17, 1.291629361630079e+17, 1.29162936166289e+17, 1.291629361695704e+17, 1.291629361726954e+17, 1.291629361759766e+17, 1.291629361791016e+17, 1.291629361823828e+17, 1.291629361856641e+17, 1.29162936188789e+17, 1.291629361920704e+17, 1.291629361951954e+17, 1.291629361984765e+17, 1.291629362017578e+17, 1.291629362048829e+17, 1.291629362081641e+17, 1.291629362114454e+17, 1.291629362145704e+17, 1.291629362178516e+17, 1.291629362209765e+17, 1.291629362242579e+17, 1.291629362275391e+17, 1.291629362306641e+17, 1.291629362339453e+17, 1.291629362370703e+17, 1.291629362403516e+17, 1.291629362436329e+17, 1.291629362467579e+17, 1.29162936250039e+17, 1.29162936253164e+17, 1.291629362564453e+17, 1.291629362597266e+17, 1.291629362628516e+17, 1.291629362661329e+17, 1.291629362694141e+17, 1.291629362725391e+17, 1.291629362758204e+17, 1.291629362789454e+17, 1.291629362822266e+17, 1.291629362855078e+17, 1.291629362886328e+17, 1.291629362919141e+17, 1.291629362950391e+17, 1.291629362983204e+17, 1.291629363014454e+17, 1.291629363047267e+17, 1.291629363080079e+17, 1.291629363111329e+17, 1.291629363144141e+17, 1.291629363176954e+17, 1.291629363208204e+17, 1.291629363241016e+17, 1.291629363272266e+17, 1.291629363305079e+17, 1.291629363336329e+17, 1.29162936336914e+17, 1.291629363401953e+17, 1.291629363433203e+17, 1.291629363466016e+17, 1.291629363498829e+17, 1.291629363530079e+17, 1.29162936356289e+17, 1.291629363594141e+17, 1.291629363626954e+17, 1.291629363658204e+17, 1.291629363691016e+17, 1.291629363723828e+17, 1.291629363755078e+17, 1.291629363787891e+17, 1.291629363819141e+17, 1.291629363851954e+17, 1.291629363884765e+17, 1.291629363916015e+17, 1.291629363948829e+17, 1.291629363981641e+17, 1.291629364012891e+17, 1.291629364045704e+17, 1.291629364076954e+17, 1.291629364109766e+17, 1.291629364142578e+17, 1.291629364173829e+17, 1.291629364206641e+17, 1.291629364237891e+17, 1.291629364270703e+17, 1.291629364303516e+17, 1.291629364334766e+17, 1.291629364367579e+17, 1.291629364398829e+17, 1.29162936443164e+17, 1.291629364464453e+17, 1.291629364495704e+17, 1.291629364528516e+17, 1.291629364559766e+17, 1.291629364592579e+17, 1.291629364625391e+17, 1.291629364656641e+17, 1.291629364689453e+17, 1.291629364722267e+17, 1.291629364753516e+17, 1.291629364786328e+17, 1.291629364817578e+17, 1.291629364850391e+17, 1.291629364883203e+17, 1.291629364914454e+17, 1.291629364947267e+17, 1.291629364978515e+17, 1.291629365011328e+17, 1.291629365044141e+17, 1.291629365075391e+17, 1.291629365108204e+17, 1.291629365139453e+17, 1.291629365172266e+17, 1.291629365205078e+17, 1.291629365236329e+17, 1.291629365269142e+17, 1.29162936530039e+17, 1.291629365333203e+17, 1.291629365366016e+17, 1.291629365397266e+17, 1.291629365430077e+17, 1.291629365461329e+17, 1.291629365494141e+17, 1.291629365526953e+17, 1.291629365558203e+17, 1.291629365591016e+17, 1.291629365622266e+17, 1.291629365655078e+17, 1.291629365687891e+17, 1.291629365719141e+17, 1.291629365751953e+17, 1.291629365783204e+17, 1.291629365816017e+17, 1.291629365848828e+17, 1.291629365880078e+17, 1.291629365912891e+17, 1.291629365944141e+17, 1.291629365976954e+17, 1.291629366009766e+17, 1.291629366041016e+17, 1.291629366073828e+17, 1.291629366105079e+17, 1.291629366137892e+17, 1.291629366170703e+17, 1.291629366201953e+17, 1.291629366234766e+17, 1.291629366267579e+17, 1.291629366298828e+17, 1.291629366331642e+17, 1.291629366362892e+17, 1.291629366395703e+17, 1.291629366426953e+17, 1.291629366459766e+17, 1.291629366492579e+17, 1.291629366523828e+17, 1.291629366556641e+17, 1.291629366589453e+17, 1.291629366620703e+17, 1.291629366653516e+17, 1.291629366684767e+17, 1.291629366717578e+17, 1.291629366748828e+17, 1.291629366781641e+17, 1.291629366814454e+17, 1.291629366845704e+17, 1.291629366878516e+17, 1.291629366909766e+17, 1.291629366942578e+17, 1.291629366975391e+17, 1.291629367006642e+17, 1.291629367039453e+17, 1.291629367070703e+17, 1.291629367103516e+17, 1.291629367136329e+17, 1.291629367167578e+17, 1.291629367200392e+17, 1.291629367231642e+17, 1.291629367264453e+17, 1.291629367297266e+17, 1.291629367328516e+17, 1.291629367361329e+17, 1.291629367392579e+17, 1.291629367425391e+17, 1.291629367458203e+17, 1.291629367489453e+17, 1.291629367522266e+17, 1.291629367555078e+17, 1.291629367586328e+17, 1.291629367619141e+17, 1.291629367650391e+17, 1.291629367683204e+17, 1.291629367714452e+17, 1.291629367747267e+17, 1.291629367780078e+17, 1.291629367811328e+17, 1.291629367844141e+17, 1.291629367876954e+17, 1.291629367908204e+17, 1.291629367941016e+17, 1.291629367972266e+17, 1.291629368005078e+17, 1.291629368036328e+17, 1.29162936806914e+17, 1.291629368101953e+17, 1.291629368133203e+17, 1.291629368166016e+17, 1.291629368198829e+17, 1.291629368230079e+17, 1.291629368262892e+17, 1.291629368295703e+17, 1.291629368326953e+17, 1.291629368359767e+17, 1.291629368391016e+17, 1.291629368423828e+17, 1.291629368455078e+17, 1.291629368487891e+17, 1.291629368520703e+17, 1.291629368551954e+17, 1.291629368584767e+17, 1.291629368616017e+17, 1.291629368648828e+17, 1.291629368681641e+17, 1.291629368712891e+17, 1.291629368745704e+17, 1.291629368776954e+17, 1.291629368809766e+17, 1.291629368842578e+17, 1.291629368873828e+17, 1.291629368906642e+17, 1.291629368937891e+17, 1.291629368970703e+17, 1.291629369003516e+17, 1.291629369034766e+17, 1.291629369067578e+17, 1.291629369100392e+17, 1.291629369131642e+17, 1.291629369164453e+17, 1.291629369195703e+17, 1.291629369228517e+17, 1.291629369261329e+17, 1.291629369292579e+17, 1.291629369325391e+17, 1.291629369356641e+17, 1.291629369389453e+17, 1.291629369422266e+17, 1.291629369453517e+17, 1.291629369486328e+17, 1.291629369517578e+17, 1.291629369550391e+17, 1.291629369583204e+17, 1.291629369614454e+17, 1.291629369647267e+17, 1.291629369678516e+17, 1.291629369711328e+17, 1.291629369744141e+17, 1.291629369775392e+17, 1.291629369808204e+17, 1.291629369839453e+17, 1.291629369872266e+17, 1.291629369905079e+17, 1.291629369936328e+17, 1.291629369969142e+17, 1.291629370000392e+17, 1.291629370033203e+17, 1.291629370066016e+17, 1.291629370097267e+17, 1.291629370130079e+17, 1.291629370161329e+17, 1.291629370194141e+17, 1.291629370226954e+17, 1.291629370258203e+17, 1.291629370291016e+17, 1.291629370322267e+17, 1.291629370355078e+17, 1.291629370387891e+17, 1.291629370419141e+17, 1.291629370451954e+17, 1.291629370483203e+17, 1.291629370516017e+17, 1.291629370548828e+17, 1.291629370580078e+17, 1.291629370612891e+17, 1.291629370644142e+17, 1.291629370676954e+17, 1.291629370709766e+17, 1.291629370741016e+17, 1.291629370773829e+17, 1.291629370805078e+17, 1.291629370837892e+17, 1.291629370870703e+17, 1.291629370901953e+17, 1.291629370934766e+17, 1.291629370966016e+17, 1.291629370998829e+17, 1.29162937103164e+17, 1.291629371062892e+17, 1.291629371095703e+17, 1.291629371128516e+17, 1.291629371159766e+17, 1.291629371192579e+17, 1.291629371223828e+17, 1.291629371256641e+17, 1.291629371289454e+17, 1.291629371320704e+17, 1.291629371353516e+17, 1.291629371384767e+17, 1.291629371417578e+17, 1.291629371448828e+17, 1.291629371481641e+17, 1.291629371514454e+17, 1.291629371545704e+17, 1.291629371578516e+17, 1.291629371611328e+17, 1.291629371642579e+17, 1.291629371675391e+17, 1.291629371706641e+17, 1.291629371739453e+17, 1.291629371772266e+17, 1.291629371803516e+17, 1.291629371836329e+17, 1.291629371867579e+17, 1.29162937190039e+17, 1.291629371933203e+17, 1.291629371964453e+17, 1.291629371997266e+17, 1.291629372028516e+17, 1.291629372061329e+17, 1.29162937209414e+17, 1.291629372125391e+17, 1.291629372158203e+17, 1.291629372189454e+17, 1.291629372222266e+17, 1.291629372255078e+17, 1.291629372286328e+17, 1.291629372319141e+17, 1.291629372350391e+17, 1.291629372383204e+17, 1.291629372416015e+17, 1.291629372447265e+17, 1.291629372480078e+17, 1.291629372511329e+17, 1.291629372544141e+17, 1.291629372576954e+17, 1.291629372608204e+17, 1.291629372641016e+17, 1.291629372672266e+17, 1.291629372705079e+17, 1.291629372737891e+17, 1.29162937276914e+17, 1.291629372801953e+17, 1.291629372834766e+17, 1.291629372866016e+17, 1.291629372898829e+17, 1.291629372930079e+17, 1.29162937296289e+17, 1.291629372995704e+17, 1.291629373026953e+17, 1.291629373059766e+17, 1.291629373091016e+17, 1.291629373123828e+17, 1.29162937315664e+17, 1.291629373187891e+17, 1.291629373220704e+17, 1.291629373251954e+17, 1.291629373284765e+17, 1.29162937331758e+17, 1.291629373348828e+17, 1.291629373381641e+17, 1.291629373412891e+17, 1.291629373445704e+17, 1.291629373478515e+17, 1.291629373509765e+17, 1.291629373542579e+17, 1.291629373573828e+17, 1.291629373606641e+17, 1.291629373639453e+17, 1.291629373670703e+17, 1.291629373703515e+17, 1.291629373734766e+17, 1.291629373767579e+17, 1.29162937380039e+17, 1.29162937383164e+17, 1.291629373864454e+17, 1.291629373895703e+17, 1.291629373928516e+17, 1.291629373961329e+17, 1.291629373992579e+17, 1.29162937402539e+17, 1.291629374056641e+17, 1.291629374089454e+17, 1.291629374122266e+17, 1.291629374153516e+17, 1.29162937418633e+17, 1.291629374217578e+17, 1.291629374250391e+17, 1.291629374283204e+17, 1.291629374314454e+17, 1.291629374347265e+17, 1.291629374378515e+17, 1.291629374411329e+17, 1.291629374444141e+17, 1.291629374475391e+17, 1.291629374508204e+17, 1.291629374541016e+17, 1.291629374572265e+17, 1.291629374605079e+17, 1.291629374636329e+17, 1.29162937466914e+17, 1.291629374701953e+17, 1.291629374733204e+17, 1.291629374766016e+17, 1.291629374798829e+17, 1.291629374830079e+17, 1.291629374862892e+17, 1.29162937489414e+17, 1.291629374926954e+17, 1.291629374959766e+17, 1.291629374991016e+17, 1.291629375023828e+17, 1.291629375056641e+17, 1.291629375087891e+17, 1.291629375120704e+17, 1.291629375151954e+17, 1.291629375184765e+17, 1.291629375216015e+17, 1.291629375248829e+17, 1.291629375281641e+17, 1.291629375312891e+17, 1.291629375345704e+17, 1.291629375376954e+17, 1.291629375409766e+17, 1.291629375442579e+17, 1.291629375473829e+17, 1.291629375506641e+17, 1.291629375539453e+17, 1.291629375570703e+17, 1.291629375603516e+17, 1.291629375634766e+17, 1.291629375667579e+17, 1.29162937570039e+17, 1.291629375731642e+17, 1.291629375764453e+17, 1.291629375795704e+17, 1.291629375828516e+17, 1.291629375861329e+17, 1.291629375892579e+17, 1.291629375925391e+17, 1.291629375956641e+17, 1.291629375989454e+17, 1.291629376022266e+17, 1.291629376053516e+17, 1.291629376086328e+17, 1.291629376117578e+17, 1.291629376150391e+17, 1.291629376183203e+17, 1.291629376214454e+17, 1.291629376247265e+17, 1.291629376278516e+17, 1.291629376311328e+17, 1.291629376344141e+17, 1.291629376375391e+17, 1.291629376408204e+17, 1.291629376439453e+17, 1.291629376472266e+17, 1.291629376505078e+17, 1.291629376536329e+17, 1.29162937656914e+17, 1.29162937660039e+17, 1.291629376633203e+17, 1.291629376664454e+17, 1.291629376697266e+17, 1.291629376730079e+17, 1.291629376761329e+17, 1.291629376794141e+17, 1.291629376826953e+17, 1.291629376858204e+17, 1.291629376891016e+17, 1.291629376923828e+17, 1.291629376955078e+17, 1.291629376987891e+17, 1.291629377019141e+17, 1.291629377051953e+17, 1.291629377083204e+17, 1.291629377116015e+17, 1.291629377148828e+17, 1.291629377180078e+17, 1.291629377212891e+17, 1.291629377244141e+17, 1.291629377276954e+17, 1.291629377309766e+17, 1.291629377341016e+17, 1.291629377373828e+17, 1.291629377405079e+17, 1.291629377437891e+17, 1.291629377470703e+17, 1.291629377501953e+17, 1.291629377534766e+17, 1.291629377566016e+17, 1.291629377598829e+17, 1.291629377631642e+17, 1.29162937766289e+17, 1.291629377695703e+17, 1.291629377726954e+17, 1.291629377759766e+17, 1.291629377792577e+17, 1.291629377823828e+17, 1.291629377856641e+17, 1.291629377887891e+17, 1.291629377920703e+17, 1.291629377953517e+17, 1.291629377984765e+17, 1.291629378017578e+17, 1.291629378048828e+17, 1.291629378081641e+17, 1.291629378114452e+17, 1.291629378145704e+17, 1.291629378178516e+17, 1.291629378211328e+17, 1.291629378242578e+17, 1.291629378275392e+17, 1.291629378306641e+17, 1.291629378339453e+17, 1.291629378372266e+17, 1.291629378403516e+17, 1.291629378436328e+17, 1.291629378469142e+17, 1.291629378500392e+17, 1.291629378533203e+17, 1.291629378564453e+17, 1.291629378597266e+17, 1.291629378630079e+17, 1.291629378661327e+17, 1.291629378694141e+17, 1.291629378725391e+17, 1.291629378758203e+17, 1.291629378789453e+17, 1.291629378822267e+17, 1.291629378855078e+17, 1.291629378886328e+17, 1.291629378919141e+17, 1.291629378951954e+17, 1.291629378983203e+17, 1.291629379016017e+17, 1.291629379047267e+17, 1.291629379080078e+17, 1.291629379112891e+17, 1.291629379144141e+17, 1.291629379176954e+17, 1.291629379208204e+17, 1.291629379241016e+17, 1.291629379273828e+17, 1.291629379305078e+17, 1.291629379337892e+17, 1.291629379369142e+17, 1.291629379401953e+17, 1.291629379434766e+17, 1.291629379466016e+17, 1.291629379498829e+17, 1.291629379531642e+17, 1.291629379562892e+17, 1.291629379595703e+17, 1.291629379626953e+17, 1.291629379659766e+17, 1.291629379692579e+17, 1.291629379723828e+17, 1.291629379756641e+17, 1.291629379787891e+17, 1.291629379820704e+17, 1.291629379853517e+17, 1.291629379884767e+17, 1.291629379917578e+17, 1.291629379948828e+17, 1.291629379981641e+17, 1.291629380014454e+17, 1.291629380045704e+17, 1.291629380078516e+17, 1.291629380109766e+17, 1.291629380142578e+17, 1.291629380173828e+17, 1.291629380206641e+17, 1.291629380239453e+17, 1.291629380270703e+17, 1.291629380303516e+17, 1.291629380336328e+17, 1.291629380367579e+17, 1.291629380400392e+17, 1.291629380431642e+17, 1.291629380464453e+17, 1.291629380495703e+17, 1.291629380528516e+17, 1.291629380561329e+17, 1.291629380592579e+17, 1.291629380625391e+17, 1.291629380656641e+17, 1.291629380689453e+17, 1.291629380722267e+17, 1.291629380753517e+17, 1.291629380786328e+17, 1.291629380817578e+17, 1.291629380850391e+17, 1.291629380883204e+17, 1.291629380914454e+17, 1.291629380947267e+17, 1.291629380978516e+17, 1.291629381011328e+17, 1.291629381044141e+17, 1.291629381075391e+17, 1.291629381108204e+17, 1.291629381139453e+17, 1.291629381172266e+17, 1.291629381205078e+17, 1.291629381236329e+17, 1.291629381269142e+17, 1.291629381300392e+17, 1.291629381333203e+17, 1.291629381366016e+17, 1.291629381397266e+17, 1.291629381430079e+17, 1.291629381461329e+17, 1.291629381494141e+17, 1.291629381526953e+17, 1.291629381558203e+17, 1.291629381591017e+17, 1.291629381622266e+17, 1.291629381655078e+17, 1.291629381687891e+17, 1.291629381719141e+17, 1.291629381751953e+17, 1.291629381783204e+17, 1.291629381816017e+17, 1.291629381848828e+17, 1.291629381880078e+17, 1.291629381912891e+17, 1.291629381945704e+17, 1.291629381976954e+17, 1.291629382009766e+17, 1.291629382041016e+17, 1.291629382073828e+17, 1.291629382105078e+17, 1.291629382137892e+17, 1.291629382170703e+17, 1.291629382201953e+17, 1.291629382234766e+17, 1.291629382266016e+17, 1.291629382298829e+17, 1.291629382331642e+17, 1.291629382362892e+17, 1.291629382395703e+17, 1.291629382426953e+17, 1.291629382459767e+17, 1.291629382492579e+17, 1.291629382523828e+17, 1.291629382556641e+17, 1.291629382587891e+17, 1.291629382620703e+17, 1.291629382653516e+17, 1.291629382684767e+17, 1.291629382717578e+17, 1.291629382750391e+17, 1.291629382781641e+17, 1.291629382814454e+17, 1.291629382845704e+17, 1.291629382878516e+17, 1.291629382911329e+17, 1.291629382942578e+17, 1.291629382975391e+17, 1.291629383006642e+17, 1.291629383039453e+17, 1.291629383072266e+17, 1.291629383103516e+17, 1.291629383136329e+17, 1.291629383167578e+17, 1.291629383200392e+17, 1.291629383233203e+17, 1.291629383264453e+17, 1.291629383297266e+17, 1.291629383328517e+17, 1.291629383361329e+17, 1.29162938339414e+17, 1.291629383425391e+17, 1.291629383458204e+17, 1.291629383489453e+17, 1.291629383522266e+17, 1.291629383555078e+17, 1.291629383586328e+17, 1.291629383619141e+17, 1.291629383650391e+17, 1.291629383683204e+17, 1.291629383716015e+17, 1.291629383747267e+17, 1.291629383780079e+17, 1.291629383811328e+17, 1.291629383844141e+17, 1.291629383876954e+17, 1.291629383908204e+17, 1.291629383941015e+17, 1.291629383972266e+17, 1.291629384005079e+17, 1.291629384037891e+17, 1.29162938406914e+17, 1.291629384101953e+17, 1.291629384133203e+17, 1.291629384166016e+17, 1.291629384198829e+17, 1.291629384230079e+17, 1.29162938426289e+17, 1.291629384294141e+17, 1.291629384326954e+17, 1.291629384359766e+17, 1.291629384391016e+17, 1.291629384423828e+17, 1.291629384455078e+17, 1.291629384487891e+17, 1.291629384520704e+17, 1.291629384551954e+17, 1.291629384584765e+17, 1.291629384616017e+17, 1.291629384648828e+17, 1.291629384681641e+17, 1.291629384712891e+17, 1.291629384745704e+17, 1.291629384776954e+17, 1.291629384809765e+17, 1.291629384842579e+17, 1.291629384873829e+17, 1.291629384906641e+17, 1.291629384937891e+17, 1.291629384970703e+17, 1.291629385003516e+17, 1.291629385034766e+17, 1.291629385067579e+17, 1.291629385098829e+17, 1.29162938513164e+17, 1.291629385164453e+17, 1.291629385195704e+17, 1.291629385228516e+17, 1.291629385259766e+17, 1.291629385292579e+17, 1.291629385325391e+17, 1.291629385356641e+17, 1.291629385389454e+17, 1.291629385420704e+17, 1.291629385453516e+17, 1.291629385486328e+17, 1.291629385517578e+17, 1.291629385550391e+17, 1.291629385581641e+17, 1.291629385614454e+17, 1.291629385647265e+17, 1.291629385678515e+17, 1.291629385711328e+17, 1.291629385744141e+17, 1.291629385775391e+17, 1.291629385808204e+17, 1.291629385839453e+17, 1.291629385872266e+17, 1.291629385905079e+17, 1.291629385936329e+17, 1.29162938596914e+17, 1.29162938600039e+17, 1.291629386033203e+17, 1.291629386066016e+17, 1.291629386097266e+17, 1.291629386130079e+17, 1.291629386161329e+17, 1.29162938619414e+17, 1.291629386226954e+17, 1.291629386258204e+17, 1.291629386291016e+17, 1.291629386322266e+17, 1.291629386355078e+17, 1.291629386387891e+17, 1.291629386419141e+17, 1.291629386451954e+17, 1.291629386483204e+17, 1.291629386516015e+17, 1.291629386548829e+17, 1.291629386580078e+17, 1.291629386612891e+17, 1.291629386644141e+17, 1.291629386676954e+17, 1.291629386709765e+17, 1.291629386741016e+17, 1.291629386773829e+17, 1.291629386805079e+17, 1.291629386837891e+17, 1.291629386870705e+17, 1.291629386901953e+17, 1.291629386934766e+17, 1.291629386967579e+17, 1.291629386998829e+17, 1.29162938703164e+17, 1.29162938706289e+17, 1.291629387095704e+17, 1.291629387128516e+17, 1.291629387159766e+17, 1.291629387192579e+17, 1.291629387223828e+17, 1.29162938725664e+17, 1.291629387289454e+17, 1.291629387320704e+17, 1.291629387353516e+17, 1.291629387384765e+17, 1.29162938741758e+17, 1.291629387450391e+17, 1.291629387481641e+17, 1.291629387514454e+17, 1.291629387545704e+17, 1.291629387578515e+17, 1.291629387611329e+17, 1.291629387642579e+17, 1.291629387675391e+17, 1.291629387706641e+17, 1.291629387739453e+17, 1.291629387772266e+17, 1.291629387803516e+17, 1.291629387836329e+17, 1.291629387867579e+17, 1.29162938790039e+17, 1.291629387933203e+17, 1.291629387964454e+17, 1.291629387997266e+17, 1.291629388028516e+17, 1.291629388061329e+17, 1.291629388094141e+17, 1.29162938812539e+17, 1.291629388158204e+17, 1.291629388189454e+17, 1.291629388222266e+17, 1.291629388255078e+17, 1.29162938828633e+17, 1.291629388319141e+17, 1.291629388350391e+17, 1.291629388383204e+17, 1.291629388416017e+17, 1.291629388447265e+17, 1.291629388480079e+17, 1.291629388511329e+17, 1.291629388544141e+17, 1.291629388576954e+17, 1.291629388608204e+17, 1.291629388641016e+17, 1.291629388672265e+17, 1.291629388705079e+17, 1.291629388737891e+17, 1.29162938876914e+17, 1.291629388801953e+17, 1.291629388833204e+17, 1.291629388866016e+17, 1.291629388898829e+17, 1.291629388930079e+17, 1.291629388962892e+17, 1.291629388995703e+17, 1.291629389026954e+17, 1.291629389059766e+17, 1.291629389091016e+17, 1.291629389123828e+17, 1.291629389156641e+17, 1.291629389187891e+17, 1.291629389220704e+17, 1.291629389251954e+17, 1.291629389284767e+17, 1.291629389317578e+17, 1.291629389348829e+17, 1.291629389381641e+17, 1.291629389412891e+17, 1.291629389445704e+17, 1.291629389478516e+17, 1.291629389509766e+17, 1.291629389542578e+17, 1.291629389575391e+17, 1.291629389606641e+17, 1.291629389639453e+17, 1.291629389670703e+17, 1.291629389703516e+17, 1.291629389736328e+17, 1.291629389767579e+17, 1.29162938980039e+17, 1.291629389831642e+17, 1.291629389864453e+17, 1.291629389897266e+17, 1.291629389928516e+17, 1.291629389961329e+17, 1.291629389994141e+17, 1.291629390025391e+17, 1.291629390058203e+17, 1.291629390089454e+17, 1.291629390122266e+17, 1.291629390155078e+17, 1.291629390186328e+17, 1.291629390219141e+17, 1.291629390250391e+17, 1.291629390283203e+17, 1.291629390314454e+17, 1.291629390347267e+17, 1.291629390380078e+17, 1.291629390411328e+17, 1.291629390444141e+17, 1.291629390476954e+17, 1.291629390508204e+17, 1.291629390541016e+17, 1.291629390572266e+17, 1.291629390605078e+17, 1.291629390636329e+17, 1.29162939066914e+17, 1.291629390701953e+17, 1.291629390733203e+17, 1.291629390766016e+17, 1.291629390798828e+17, 1.291629390830079e+17, 1.291629390862892e+17, 1.291629390894141e+17, 1.291629390926953e+17, 1.291629390959767e+17, 1.291629390991016e+17, 1.291629391023828e+17, 1.291629391055078e+17, 1.291629391087891e+17, 1.291629391119141e+17, 1.291629391151953e+17, 1.291629391184767e+17, 1.291629391216015e+17, 1.291629391248828e+17, 1.291629391280078e+17, 1.291629391312891e+17, 1.291629391345702e+17, 1.291629391376954e+17, 1.291629391409766e+17, 1.291629391441016e+17, 1.291629391473828e+17, 1.291629391506642e+17, 1.291629391537891e+17, 1.291629391570703e+17, 1.291629391601953e+17, 1.291629391634766e+17, 1.291629391667578e+17, 1.291629391698828e+17, 1.291629391731642e+17, 1.291629391764453e+17, 1.291629391795703e+17, 1.291629391828516e+17, 1.291629391859766e+17, 1.291629391892579e+17, 1.291629391925391e+17, 1.291629391956641e+17, 1.291629391989453e+17, 1.291629392022267e+17, 1.291629392053517e+17, 1.291629392086328e+17, 1.291629392117578e+17, 1.291629392150391e+17, 1.291629392183204e+17, 1.291629392214452e+17, 1.291629392247267e+17, 1.291629392280078e+17, 1.291629392311328e+17, 1.291629392344141e+17, 1.291629392375392e+17, 1.291629392408204e+17, 1.291629392439453e+17, 1.291629392472266e+17, 1.291629392505079e+17, 1.291629392536328e+17, 1.291629392569142e+17, 1.291629392601953e+17, 1.291629392633203e+17, 1.291629392666016e+17, 1.291629392697266e+17, 1.291629392730079e+17, 1.291629392762892e+17, 1.291629392794141e+17, 1.291629392826953e+17, 1.291629392858203e+17, 1.291629392891016e+17, 1.291629392923828e+17, 1.291629392955078e+17, 1.291629392987891e+17, 1.291629393019141e+17, 1.291629393051954e+17, 1.291629393084767e+17, 1.291629393116017e+17, 1.291629393148828e+17, 1.291629393180078e+17, 1.291629393212891e+17, 1.291629393245704e+17, 1.291629393276954e+17, 1.291629393309766e+17, 1.291629393342578e+17, 1.291629393373829e+17, 1.291629393406641e+17, 1.291629393437892e+17, 1.291629393470703e+17, 1.291629393503516e+17, 1.291629393534766e+17, 1.291629393567579e+17, 1.291629393598829e+17, 1.291629393631642e+17, 1.291629393664453e+17, 1.291629393695703e+17, 1.291629393728516e+17, 1.291629393759766e+17, 1.291629393792579e+17, 1.291629393825391e+17, 1.291629393856641e+17, 1.291629393889453e+17, 1.291629393920704e+17, 1.291629393953517e+17, 1.291629393986328e+17, 1.291629394017578e+17, 1.291629394050391e+17, 1.291629394081641e+17, 1.291629394114454e+17, 1.291629394145704e+17, 1.291629394178516e+17, 1.291629394211328e+17, 1.291629394242578e+17, 1.291629394275391e+17, 1.291629394306641e+17, 1.291629394339453e+17, 1.291629394372266e+17, 1.291629394403516e+17, 1.291629394436328e+17, 1.291629394467579e+17, 1.291629394500392e+17, 1.291629394533203e+17, 1.291629394564453e+17, 1.291629394597266e+17, 1.291629394628516e+17, 1.291629394661329e+17, 1.291629394692579e+17, 1.291629394725391e+17, 1.291629394758203e+17, 1.291629394789454e+17, 1.291629394822267e+17, 1.291629394853517e+17, 1.291629394886328e+17, 1.291629394919141e+17, 1.291629394950391e+17, 1.291629394983204e+17, 1.291629395014454e+17, 1.291629395047267e+17, 1.291629395080078e+17, 1.291629395111328e+17, 1.291629395144141e+17, 1.291629395176954e+17, 1.291629395208204e+17, 1.291629395241016e+17, 1.291629395272266e+17, 1.291629395305078e+17, 1.291629395336329e+17, 1.291629395369142e+17, 1.291629395401953e+17, 1.291629395434766e+17, 1.291629395466016e+17, 1.291629395498829e+17, 1.29162939553164e+17, 1.291629395564453e+17, 1.291629395597266e+17, 1.291629395628516e+17, 1.291629395661329e+17, 1.29162939569414e+17, 1.291629395726953e+17, 1.291629395759766e+17, 1.291629395791016e+17, 1.291629395823828e+17, 1.291629395858203e+17, 1.291629395891016e+17, 1.291629395922267e+17, 1.291629395955078e+17, 1.291629395986328e+17, 1.291629396019141e+17, 1.291629396051954e+17, 1.291629396084765e+17, 1.291629396116017e+17, 1.291629396148828e+17, 1.291629396181641e+17, 1.291629396214454e+17, 1.291629396247265e+17, 1.291629396278515e+17, 1.291629396311329e+17, 1.291629396344141e+17, 1.291629396375391e+17, 1.291629396408204e+17, 1.291629396439453e+17, 1.291629396472266e+17, 1.291629396505079e+17, 1.291629396536329e+17, 1.29162939656914e+17, 1.291629396601953e+17, 1.291629396633204e+17, 1.291629396666016e+17, 1.291629396697266e+17, 1.291629396730079e+17, 1.291629396762892e+17, 1.29162939679414e+17, 1.291629396826954e+17, 1.291629396858204e+17, 1.291629396891016e+17, 1.291629396923828e+17, 1.29162939695508e+17, 1.291629396987891e+17, 1.291629397019141e+17, 1.291629397051954e+17, 1.291629397084767e+17, 1.291629397116015e+17, 1.291629397148828e+17, 1.291629397181641e+17, 1.291629397212891e+17, 1.291629397245704e+17, 1.291629397276954e+17, 1.291629397309766e+17, 1.291629397342578e+17, 1.291629397373829e+17, 1.291629397406641e+17, 1.291629397437891e+17, 1.291629397470703e+17, 1.291629397503516e+17, 1.291629397534766e+17, 1.291629397567579e+17, 1.291629397598829e+17, 1.291629397631642e+17, 1.291629397664453e+17, 1.291629397695704e+17, 1.291629397728516e+17, 1.291629397759766e+17, 1.291629397792579e+17, 1.29162939782383e+17, 1.291629397856641e+17, 1.291629397889453e+17, 1.291629397920704e+17, 1.291629397953517e+17, 1.291629397986328e+17, 1.291629398017578e+17, 1.291629398050391e+17, 1.291629398081641e+17, 1.291629398114454e+17, 1.291629398147267e+17, 1.291629398178516e+17, 1.291629398211328e+17, 1.291629398242579e+17, 1.291629398275391e+17, 1.291629398308204e+17, 1.291629398339453e+17, 1.291629398372266e+17, 1.291629398403516e+17, 1.291629398436329e+17, 1.29162939846914e+17, 1.291629398500392e+17, 1.291629398533203e+17, 1.291629398564453e+17, 1.291629398597266e+17, 1.291629398630079e+17, 1.291629398661329e+17, 1.291629398694141e+17, 1.291629398725391e+17, 1.291629398758203e+17, 1.291629398791016e+17, 1.291629398822266e+17, 1.291629398855078e+17, 1.291629398886328e+17, 1.291629398919141e+17, 1.291629398951953e+17, 1.291629398983204e+17, 1.291629399016015e+17, 1.291629399047267e+17, 1.291629399080078e+17, 1.291629399112891e+17, 1.291629399144141e+17, 1.291629399176954e+17, 1.291629399208204e+17, 1.291629399241016e+17, 1.291629399273828e+17, 1.291629399305078e+17, 1.291629399337891e+17, 1.291629399369142e+17, 1.291629399401953e+17, 1.291629399434766e+17, 1.291629399466016e+17, 1.291629399498829e+17, 1.291629399530079e+17, 1.291629399562892e+17, 1.291629399595703e+17, 1.291629399626953e+17, 1.291629399659766e+17, 1.291629399691016e+17, 1.291629399723828e+17, 1.291629399756641e+17, 1.291629399787891e+17, 1.291629399820703e+17, 1.291629399851954e+17, 1.291629399884765e+17, 1.291629399917578e+17, 1.291629399948828e+17, 1.291629399981641e+17, 1.291629400012891e+17, 1.291629400045704e+17, 1.291629400078516e+17, 1.291629400109766e+17, 1.291629400142578e+17, 1.291629400173828e+17, 1.291629400206641e+17, 1.291629400239453e+17, 1.291629400270703e+17, 1.291629400303516e+17, 1.291629400336328e+17, 1.291629400367578e+17, 1.291629400400392e+17, 1.291629400431642e+17, 1.291629400464453e+17, 1.291629400495703e+17, 1.291629400528516e+17, 1.291629400561329e+17, 1.291629400592579e+17, 1.291629400625391e+17, 1.291629400656641e+17, 1.291629400689453e+17, 1.291629400722267e+17, 1.291629400753516e+17, 1.291629400786328e+17, 1.291629400819141e+17, 1.291629400850391e+17, 1.291629400883203e+17, 1.291629400914454e+17, 1.291629400947267e+17, 1.291629400980078e+17, 1.291629401011328e+17, 1.291629401044142e+17, 1.291629401075391e+17, 1.291629401108204e+17, 1.291629401141016e+17, 1.291629401172266e+17, 1.291629401205078e+17, 1.291629401236328e+17, 1.291629401269142e+17, 1.291629401301953e+17, 1.291629401333203e+17, 1.291629401366016e+17, 1.291629401397266e+17, 1.291629401430077e+17, 1.291629401462892e+17, 1.291629401494141e+17, 1.291629401526953e+17, 1.291629401558203e+17, 1.291629401591017e+17, 1.291629401623828e+17, 1.291629401655078e+17, 1.291629401687891e+17, 1.291629401719141e+17, 1.291629401751953e+17, 1.291629401783203e+17, 1.291629401816017e+17, 1.291629401848828e+17, 1.291629401880078e+17, 1.291629401912891e+17, 1.291629401945704e+17, 1.291629401976954e+17, 1.291629402009766e+17, 1.291629402041016e+17, 1.291629402073828e+17, 1.291629402106642e+17, 1.291629402137892e+17, 1.291629402170703e+17, 1.291629402201953e+17, 1.291629402234766e+17, 1.291629402267579e+17, 1.291629402298828e+17, 1.291629402331642e+17, 1.291629402362892e+17, 1.291629402395703e+17, 1.291629402426953e+17, 1.291629402459767e+17, 1.291629402492579e+17, 1.291629402523828e+17, 1.291629402556641e+17, 1.291629402587891e+17, 1.291629402620703e+17, 1.291629402653517e+17, 1.291629402684767e+17, 1.291629402717578e+17, 1.291629402748828e+17, 1.291629402781641e+17, 1.291629402814454e+17, 1.291629402845702e+17, 1.291629402878516e+17, 1.291629402909766e+17, 1.291629402942578e+17, 1.291629402973828e+17, 1.291629403006642e+17, 1.291629403039453e+17, 1.291629403072266e+17, 1.291629403103516e+17, 1.291629403136329e+17, 1.291629403167578e+17, 1.291629403200392e+17, 1.291629403233203e+17, 1.291629403264453e+17, 1.291629403297266e+17, 1.291629403328517e+17, 1.291629403361329e+17, 1.291629403394141e+17, 1.291629403425391e+17, 1.291629403458204e+17, 1.291629403489453e+17, 1.291629403522267e+17, 1.291629403555078e+17, 1.291629403586328e+17, 1.291629403619141e+17, 1.291629403650391e+17, 1.291629403683204e+17, 1.291629403716017e+17, 1.291629403747267e+17, 1.291629403780078e+17, 1.291629403811328e+17, 1.291629403844141e+17, 1.291629403876954e+17, 1.291629403908204e+17, 1.291629403941016e+17, 1.291629403972266e+17, 1.291629404005079e+17, 1.291629404037891e+17, 1.291629404069142e+17, 1.291629404101953e+17, 1.291629404134766e+17, 1.291629404166016e+17, 1.291629404198829e+17, 1.291629404230079e+17, 1.291629404262892e+17, 1.291629404295703e+17, 1.291629404326953e+17, 1.291629404359766e+17, 1.291629404391016e+17, 1.291629404423828e+17, 1.291629404456641e+17, 1.291629404487891e+17, 1.291629404520703e+17, 1.291629404551954e+17, 1.291629404584767e+17, 1.291629404617578e+17, 1.291629404648828e+17, 1.291629404681641e+17, 1.291629404712891e+17, 1.291629404745704e+17, 1.291629404778515e+17, 1.291629404809766e+17, 1.291629404842578e+17, 1.291629404873829e+17, 1.291629404906641e+17, 1.291629404939453e+17, 1.291629404970703e+17, 1.291629405003516e+17, 1.291629405034766e+17, 1.291629405067579e+17, 1.291629405098829e+17, 1.291629405131642e+17, 1.291629405164453e+17, 1.291629405195703e+17, 1.291629405228516e+17, 1.291629405261329e+17, 1.291629405292579e+17, 1.291629405325391e+17, 1.291629405356641e+17, 1.291629405389453e+17, 1.291629405422266e+17, 1.291629405453517e+17, 1.291629405486328e+17, 1.291629405517578e+17, 1.291629405550391e+17, 1.291629405583204e+17, 1.291629405614454e+17, 1.291629405647265e+17, 1.291629405678516e+17, 1.291629405711328e+17, 1.291629405744141e+17, 1.291629405775391e+17, 1.291629405808204e+17, 1.291629405839453e+17, 1.291629405872266e+17, 1.291629405905079e+17, 1.291629405936329e+17, 1.29162940596914e+17, 1.291629406000392e+17, 1.291629406033203e+17, 1.291629406066016e+17, 1.291629406097266e+17, 1.291629406130079e+17, 1.291629406161329e+17, 1.29162940619414e+17, 1.291629406226954e+17, 1.291629406258203e+17, 1.291629406291016e+17, 1.291629406322266e+17, 1.291629406355078e+17, 1.291629406386328e+17, 1.291629406419141e+17, 1.291629406451954e+17, 1.291629406483204e+17, 1.291629406516015e+17, 1.291629406548829e+17, 1.291629406581641e+17, 1.291629406612891e+17, 1.291629406645704e+17, 1.291629406676954e+17, 1.291629406709765e+17, 1.291629406742579e+17, 1.291629406773829e+17, 1.291629406806641e+17, 1.291629406837891e+17, 1.291629406870703e+17, 1.291629406903516e+17, 1.291629406934765e+17, 1.291629406967579e+17, 1.291629406998829e+17, 1.29162940703164e+17, 1.291629407064453e+17, 1.291629407095704e+17, 1.291629407128516e+17, 1.291629407159766e+17, 1.291629407192579e+17, 1.291629407223828e+17, 1.29162940725664e+17, 1.291629407289454e+17, 1.291629407320704e+17, 1.291629407353516e+17, 1.291629407386328e+17, 1.291629407417578e+17, 1.291629407450391e+17, 1.291629407481641e+17, 1.291629407514454e+17, 1.291629407547267e+17, 1.291629407578515e+17, 1.291629407611329e+17, 1.291629407644141e+17, 1.291629407675391e+17, 1.291629407708204e+17, 1.291629407739453e+17, 1.291629407772266e+17, 1.291629407803515e+17, 1.291629407836329e+17, 1.29162940786914e+17, 1.29162940790039e+17, 1.291629407933203e+17, 1.291629407966016e+17, 1.291629407997266e+17, 1.291629408030079e+17, 1.291629408061329e+17, 1.291629408094141e+17, 1.291629408126954e+17, 1.291629408158204e+17, 1.291629408191016e+17, 1.291629408222266e+17, 1.291629408255078e+17, 1.291629408287891e+17, 1.291629408319141e+17, 1.291629408351954e+17, 1.291629408383204e+17, 1.291629408416015e+17, 1.291629408448829e+17, 1.291629408480078e+17, 1.291629408512891e+17, 1.291629408544141e+17, 1.291629408576954e+17, 1.291629408609765e+17, 1.291629408641016e+17, 1.291629408673829e+17, 1.291629408705079e+17, 1.291629408737891e+17, 1.291629408770703e+17, 1.291629408801953e+17, 1.291629408834766e+17, 1.291629408866016e+17, 1.291629408898829e+17, 1.29162940893164e+17, 1.291629408962892e+17, 1.291629408995704e+17, 1.291629409026954e+17, 1.291629409059766e+17, 1.291629409092579e+17, 1.291629409123828e+17, 1.291629409156641e+17, 1.291629409189454e+17, 1.291629409220704e+17, 1.291629409253516e+17, 1.291629409284765e+17, 1.29162940931758e+17, 1.291629409348828e+17, 1.291629409381641e+17, 1.291629409414454e+17, 1.291629409445704e+17, 1.291629409478515e+17, 1.291629409509766e+17, 1.291629409542579e+17, 1.291629409575391e+17, 1.291629409606641e+17, 1.291629409639453e+17, 1.291629409670703e+17, 1.291629409703516e+17, 1.291629409736329e+17, 1.291629409767579e+17, 1.29162940980039e+17, 1.29162940983164e+17, 1.291629409864454e+17, 1.291629409897266e+17, 1.291629409928516e+17, 1.291629409961329e+17, 1.291629409994141e+17, 1.29162941002539e+17, 1.291629410058204e+17, 1.291629410089454e+17, 1.291629410122266e+17, 1.291629410155078e+17, 1.29162941018633e+17, 1.291629410219141e+17, 1.291629410250391e+17, 1.291629410283204e+17, 1.291629410314454e+17, 1.291629410347265e+17, 1.291629410380078e+17, 1.291629410411329e+17, 1.291629410444141e+17, 1.291629410476954e+17, 1.291629410508204e+17, 1.291629410541016e+17, 1.291629410572266e+17, 1.291629410605079e+17, 1.291629410637892e+17, 1.29162941066914e+17, 1.291629410701953e+17, 1.291629410733204e+17, 1.291629410766016e+17, 1.291629410798828e+17, 1.291629410830079e+17, 1.291629410862892e+17, 1.29162941089414e+17, 1.291629410926953e+17, 1.291629410959766e+17, 1.291629410991016e+17, 1.291629411023828e+17, 1.291629411055078e+17, 1.291629411087891e+17, 1.291629411120703e+17, 1.291629411151954e+17, 1.291629411184767e+17, 1.291629411216015e+17, 1.291629411248828e+17, 1.291629411281641e+17, 1.291629411312891e+17, 1.291629411345704e+17, 1.291629411376954e+17, 1.291629411409766e+17, 1.291629411442578e+17, 1.291629411473829e+17, 1.291629411506641e+17, 1.291629411537891e+17, 1.291629411570703e+17, 1.291629411603516e+17, 1.291629411634766e+17, 1.291629411667578e+17, 1.291629411698829e+17, 1.291629411731642e+17, 1.291629411764453e+17, 1.291629411795703e+17, 1.291629411828516e+17, 1.291629411861329e+17, 1.291629411892579e+17, 1.291629411925391e+17, 1.291629411956641e+17, 1.291629411989453e+17, 1.291629412022266e+17, 1.291629412053517e+17, 1.291629412086328e+17, 1.291629412117578e+17, 1.291629412150391e+17, 1.291629412183204e+17, 1.291629412214454e+17, 1.291629412247267e+17, 1.291629412280078e+17, 1.291629412311328e+17, 1.291629412344141e+17, 1.291629412375391e+17, 1.291629412408204e+17, 1.291629412439453e+17, 1.291629412472266e+17, 1.291629412505078e+17, 1.291629412536328e+17, 1.29162941256914e+17, 1.291629412601953e+17, 1.291629412633203e+17, 1.291629412666016e+17, 1.291629412697266e+17, 1.291629412730079e+17, 1.291629412761329e+17, 1.291629412794141e+17, 1.291629412826953e+17, 1.291629412858203e+17, 1.291629412891016e+17, 1.291629412923828e+17, 1.291629412955078e+17, 1.291629412987891e+17, 1.291629413020703e+17, 1.291629413051953e+17, 1.291629413084767e+17, 1.291629413116017e+17, 1.291629413148828e+17, 1.291629413181642e+17, 1.291629413212891e+17, 1.291629413245704e+17, 1.291629413276954e+17, 1.291629413309766e+17, 1.291629413341016e+17, 1.291629413373828e+17, 1.291629413406642e+17, 1.291629413437891e+17, 1.291629413470703e+17, 1.291629413501953e+17, 1.291629413534766e+17, 1.291629413567578e+17, 1.291629413598829e+17, 1.291629413631642e+17, 1.291629413662892e+17, 1.291629413695703e+17, 1.291629413728517e+17, 1.291629413759766e+17, 1.291629413792579e+17, 1.291629413823828e+17, 1.291629413856641e+17, 1.291629413889453e+17, 1.291629413920703e+17, 1.291629413953517e+17, 1.291629413984765e+17, 1.291629414017578e+17, 1.291629414050391e+17, 1.291629414081641e+17, 1.291629414114452e+17, 1.291629414145704e+17, 1.291629414178516e+17, 1.291629414211328e+17, 1.291629414242578e+17, 1.291629414275392e+17, 1.291629414306641e+17, 1.291629414339453e+17, 1.291629414372266e+17, 1.291629414403516e+17, 1.291629414436328e+17, 1.291629414467579e+17, 1.291629414500392e+17, 1.291629414533203e+17, 1.291629414564453e+17, 1.291629414597267e+17, 1.291629414628516e+17, 1.291629414661329e+17, 1.291629414694141e+17, 1.291629414725391e+17, 1.291629414758203e+17, 1.291629414789453e+17, 1.291629414822267e+17, 1.291629414855078e+17, 1.291629414886328e+17, 1.291629414919141e+17, 1.291629414950391e+17, 1.291629414983203e+17, 1.291629415016017e+17, 1.291629415047267e+17, 1.291629415080078e+17, 1.291629415111328e+17, 1.291629415144142e+17, 1.291629415176954e+17, 1.291629415208204e+17, 1.291629415241016e+17, 1.291629415272266e+17, 1.291629415305078e+17, 1.291629415336328e+17, 1.291629415369142e+17, 1.291629415401953e+17, 1.291629415433203e+17, 1.291629415466016e+17, 1.291629415498829e+17, 1.291629415530077e+17, 1.291629415562892e+17, 1.291629415594141e+17, 1.291629415626953e+17, 1.291629415659766e+17, 1.291629415691017e+17, 1.291629415723828e+17, 1.291629415755078e+17, 1.291629415787891e+17, 1.291629415819141e+17, 1.291629415851953e+17, 1.291629415884767e+17, 1.291629415916017e+17, 1.291629415948828e+17, 1.291629415980078e+17, 1.291629416012892e+17, 1.291629416045704e+17, 1.291629416076954e+17, 1.291629416109766e+17, 1.291629416141016e+17, 1.291629416173828e+17, 1.291629416206642e+17, 1.291629416237892e+17, 1.291629416270703e+17, 1.291629416301953e+17, 1.291629416334766e+17, 1.291629416367579e+17, 1.291629416398828e+17, 1.291629416431642e+17, 1.291629416464453e+17, 1.291629416495703e+17, 1.291629416528516e+17, 1.291629416559767e+17, 1.291629416592579e+17, 1.291629416625391e+17, 1.291629416656641e+17, 1.291629416689454e+17, 1.291629416720703e+17, 1.291629416753517e+17, 1.291629416786328e+17, 1.291629416817578e+17, 1.291629416850391e+17, 1.291629416881641e+17, 1.291629416914454e+17, 1.291629416947267e+17, 1.291629416978516e+17, 1.291629417011328e+17, 1.291629417042578e+17, 1.291629417075392e+17, 1.291629417108204e+17, 1.291629417139453e+17, 1.291629417172266e+17, 1.291629417203516e+17, 1.291629417236329e+17, 1.29162941726914e+17, 1.291629417300392e+17, 1.291629417333203e+17, 1.291629417366016e+17, 1.291629417397266e+17, 1.291629417430079e+17, 1.291629417461329e+17, 1.291629417494141e+17, 1.291629417526953e+17, 1.291629417558204e+17, 1.291629417591016e+17, 1.291629417622267e+17, 1.291629417655078e+17, 1.291629417687891e+17, 1.291629417719141e+17, 1.291629417751954e+17, 1.291629417783204e+17, 1.291629417816017e+17, 1.291629417848828e+17, 1.291629417880078e+17, 1.291629417912891e+17, 1.291629417944141e+17, 1.291629417976954e+17, 1.291629418009765e+17, 1.291629418041016e+17, 1.291629418073828e+17, 1.291629418106641e+17, 1.291629418137891e+17, 1.291629418170703e+17, 1.291629418201953e+17, 1.291629418234766e+17, 1.291629418267579e+17, 1.291629418298829e+17, 1.29162941833164e+17, 1.291629418362892e+17, 1.291629418395703e+17, 1.291629418428516e+17, 1.291629418459766e+17, 1.291629418492579e+17, 1.291629418523828e+17, 1.29162941855664e+17, 1.291629418589454e+17, 1.291629418620704e+17, 1.291629418653516e+17, 1.291629418684765e+17, 1.291629418717578e+17, 1.291629418750391e+17, 1.291629418781641e+17, 1.291629418814454e+17, 1.291629418845704e+17, 1.291629418878515e+17, 1.291629418911329e+17, 1.291629418942578e+17, 1.291629418975391e+17, 1.291629419006641e+17, 1.291629419039453e+17, 1.291629419072265e+17, 1.291629419103516e+17, 1.291629419136329e+17, 1.291629419167579e+17, 1.29162941920039e+17, 1.291629419233204e+17, 1.291629419264453e+17, 1.291629419297266e+17, 1.291629419328516e+17, 1.291629419361329e+17, 1.29162941939414e+17, 1.29162941942539e+17, 1.291629419458204e+17, 1.291629419489453e+17, 1.291629419522266e+17, 1.291629419555078e+17, 1.291629419586328e+17, 1.29162941961914e+17, 1.291629419650391e+17, 1.291629419683204e+17, 1.291629419716015e+17, 1.291629419747265e+17, 1.291629419780079e+17, 1.291629419811328e+17, 1.291629419844141e+17, 1.291629419876954e+17, 1.291629419908204e+17, 1.291629419941015e+17, 1.291629419972266e+17, 1.291629420005079e+17, 1.291629420037891e+17, 1.29162942006914e+17, 1.291629420101955e+17, 1.291629420134766e+17, 1.291629420166016e+17, 1.291629420198829e+17, 1.291629420230079e+17, 1.29162942026289e+17, 1.291629420295704e+17, 1.291629420326954e+17, 1.291629420359766e+17, 1.291629420391016e+17, 1.291629420423828e+17, 1.291629420456641e+17, 1.29162942048789e+17, 1.291629420520704e+17, 1.291629420551954e+17, 1.291629420584765e+17, 1.291629420617578e+17, 1.291629420648829e+17, 1.291629420681641e+17, 1.291629420712891e+17, 1.291629420745704e+17, 1.291629420778516e+17, 1.291629420809765e+17, 1.291629420842579e+17, 1.291629420873829e+17, 1.291629420906641e+17, 1.291629420939453e+17, 1.291629420970703e+17, 1.291629421003516e+17, 1.291629421034765e+17, 1.291629421067579e+17, 1.29162942110039e+17, 1.29162942113164e+17, 1.291629421164453e+17, 1.291629421195704e+17, 1.291629421228516e+17, 1.291629421261329e+17, 1.291629421292579e+17, 1.291629421325391e+17, 1.29162942135664e+17, 1.291629421389454e+17, 1.291629421422266e+17, 1.291629421453516e+17, 1.291629421486328e+17, 1.29162942151758e+17, 1.291629421550391e+17, 1.291629421583204e+17, 1.291629421614454e+17, 1.291629421647267e+17, 1.291629421678515e+17, 1.291629421711329e+17, 1.291629421744141e+17, 1.291629421775391e+17, 1.291629421808204e+17, 1.291629421841016e+17, 1.291629421872266e+17, 1.291629421905079e+17, 1.291629421936329e+17, 1.29162942196914e+17, 1.291629422001953e+17, 1.291629422033203e+17, 1.291629422066016e+17, 1.291629422097266e+17, 1.291629422130079e+17, 1.29162942216289e+17, 1.291629422194141e+17, 1.291629422226954e+17, 1.291629422258204e+17, 1.291629422291016e+17, 1.291629422323828e+17, 1.291629422355078e+17, 1.291629422387891e+17, 1.291629422419141e+17, 1.291629422451954e+17, 1.291629422484765e+17, 1.291629422516015e+17, 1.291629422548828e+17, 1.291629422580079e+17, 1.291629422612891e+17, 1.291629422645704e+17, 1.291629422676954e+17, 1.291629422709766e+17, 1.291629422741016e+17, 1.291629422773829e+17, 1.291629422806641e+17, 1.291629422837891e+17, 1.291629422870703e+17, 1.291629422901953e+17, 1.291629422934766e+17, 1.291629422967579e+17, 1.291629422998829e+17, 1.29162942303164e+17, 1.291629423062892e+17, 1.291629423095704e+17, 1.291629423128516e+17, 1.291629423159766e+17, 1.291629423192579e+17, 1.291629423223828e+17, 1.291629423256641e+17, 1.291629423289453e+17, 1.291629423320704e+17, 1.291629423353516e+17, 1.291629423384765e+17, 1.291629423417578e+17, 1.291629423448828e+17, 1.291629423481641e+17, 1.291629423514454e+17, 1.291629423547267e+17, 1.291629423578515e+17, 1.291629423611328e+17, 1.291629423642579e+17, 1.291629423675391e+17, 1.291629423708204e+17, 1.291629423739453e+17, 1.291629423772266e+17, 1.291629423803516e+17, 1.291629423836329e+17, 1.291629423869142e+17, 1.29162942390039e+17, 1.291629423933203e+17, 1.291629423964454e+17, 1.291629423997266e+17, 1.291629424030077e+17, 1.291629424061329e+17, 1.291629424094141e+17, 1.291629424126953e+17, 1.291629424158203e+17, 1.291629424191017e+17, 1.291629424222266e+17, 1.291629424255078e+17, 1.291629424287891e+17, 1.291629424319141e+17, 1.291629424351953e+17, 1.291629424383204e+17, 1.291629424416017e+17, 1.291629424448828e+17, 1.291629424480078e+17, 1.291629424512891e+17, 1.291629424544141e+17, 1.291629424576954e+17, 1.291629424609766e+17, 1.291629424641016e+17, 1.291629424673828e+17, 1.291629424705079e+17, 1.291629424737892e+17, 1.291629424770703e+17, 1.291629424801953e+17, 1.291629424834766e+17, 1.291629424866016e+17, 1.291629424898828e+17, 1.291629424931642e+17, 1.291629424962892e+17, 1.291629424995703e+17, 1.291629425026953e+17, 1.291629425059766e+17, 1.291629425092579e+17, 1.291629425123828e+17, 1.291629425156641e+17, 1.291629425187891e+17, 1.291629425220703e+17, 1.291629425253516e+17, 1.291629425284767e+17, 1.291629425317578e+17, 1.291629425348828e+17, 1.291629425381641e+17, 1.291629425414454e+17, 1.291629425445704e+17, 1.291629425478516e+17, 1.291629425509766e+17, 1.291629425542578e+17, 1.291629425575391e+17, 1.291629425606642e+17, 1.291629425639453e+17, 1.291629425670703e+17, 1.291629425703516e+17, 1.291629425736329e+17, 1.291629425767578e+17, 1.291629425800392e+17, 1.291629425833203e+17, 1.291629425864453e+17, 1.291629425897266e+17, 1.291629425928516e+17, 1.291629425961329e+17, 1.291629425994141e+17, 1.291629426025391e+17, 1.291629426058203e+17, 1.291629426089453e+17, 1.291629426122266e+17, 1.291629426155078e+17, 1.291629426186328e+17, 1.291629426219141e+17, 1.291629426251953e+17, 1.291629426283204e+17, 1.291629426316017e+17, 1.291629426347267e+17, 1.291629426380078e+17, 1.291629426412892e+17, 1.291629426444141e+17, 1.291629426476954e+17, 1.291629426508204e+17, 1.291629426541016e+17, 1.291629426573828e+17, 1.291629426605078e+17, 1.291629426637892e+17, 1.29162942666914e+17, 1.291629426701953e+17, 1.291629426734766e+17, 1.291629426766016e+17, 1.291629426798829e+17, 1.291629426830079e+17, 1.291629426862892e+17, 1.291629426895703e+17, 1.291629426926953e+17, 1.291629426959767e+17, 1.291629426991016e+17, 1.291629427023828e+17, 1.291629427056641e+17, 1.291629427087891e+17, 1.291629427120703e+17, 1.291629427151954e+17, 1.291629427184767e+17, 1.291629427217578e+17, 1.291629427248828e+17, 1.291629427281641e+17, 1.291629427312891e+17, 1.291629427345704e+17, 1.291629427378516e+17, 1.291629427409766e+17, 1.291629427442578e+17, 1.291629427473828e+17, 1.291629427506642e+17, 1.291629427539453e+17, 1.291629427570703e+17, 1.291629427603516e+17, 1.291629427634766e+17, 1.291629427667578e+17, 1.291629427700392e+17, 1.291629427731642e+17, 1.291629427764453e+17, 1.291629427795703e+17, 1.291629427828517e+17, 1.291629427861329e+17, 1.291629427892579e+17, 1.291629427925391e+17, 1.291629427956641e+17, 1.291629427989453e+17, 1.291629428022266e+17, 1.291629428053517e+17, 1.291629428086328e+17, 1.291629428117578e+17, 1.291629428150391e+17, 1.291629428183204e+17, 1.291629428214454e+17, 1.291629428247267e+17, 1.291629428278516e+17, 1.291629428311328e+17, 1.291629428344141e+17, 1.291629428375392e+17, 1.291629428408204e+17, 1.291629428439453e+17, 1.291629428472266e+17, 1.291629428505079e+17, 1.291629428536328e+17, 1.291629428569142e+17, 1.291629428600392e+17, 1.291629428633203e+17, 1.291629428666016e+17, 1.291629428697267e+17, 1.291629428730079e+17, 1.291629428761329e+17, 1.291629428794141e+17, 1.291629428826954e+17, 1.291629428858203e+17, 1.291629428891016e+17, 1.291629428922267e+17, 1.291629428955078e+17, 1.291629428987891e+17, 1.291629429019141e+17, 1.291629429051954e+17, 1.291629429083203e+17, 1.291629429116017e+17, 1.291629429148828e+17, 1.291629429180078e+17, 1.291629429212891e+17, 1.291629429244142e+17, 1.291629429276954e+17, 1.291629429309766e+17, 1.291629429341016e+17, 1.291629429373829e+17, 1.291629429405078e+17, 1.291629429437892e+17, 1.291629429470703e+17, 1.291629429501953e+17, 1.291629429534766e+17, 1.291629429566016e+17, 1.291629429598829e+17, 1.29162942963164e+17, 1.291629429662892e+17, 1.291629429695704e+17, 1.291629429726953e+17, 1.291629429759766e+17, 1.291629429792579e+17, 1.291629429823828e+17, 1.291629429856641e+17, 1.291629429887891e+17, 1.291629429920704e+17, 1.291629429953516e+17, 1.291629429984767e+17, 1.291629430017578e+17, 1.291629430048828e+17, 1.291629430081641e+17, 1.291629430114454e+17, 1.291629430145704e+17, 1.291629430178515e+17, 1.291629430209766e+17, 1.291629430242579e+17, 1.291629430275391e+17, 1.291629430306641e+17, 1.291629430339453e+17, 1.291629430372266e+17, 1.291629430403516e+17, 1.291629430436329e+17, 1.291629430467579e+17, 1.29162943050039e+17, 1.291629430533203e+17, 1.291629430564453e+17, 1.291629430597266e+17, 1.291629430630079e+17, 1.291629430661329e+17, 1.29162943069414e+17, 1.291629430725391e+17, 1.291629430758203e+17, 1.291629430789454e+17, 1.291629430822266e+17, 1.291629430855078e+17, 1.291629430886328e+17, 1.291629430919141e+17, 1.291629430950391e+17, 1.291629430983204e+17, 1.291629431016015e+17, 1.291629431047265e+17, 1.291629431080078e+17, 1.291629431111329e+17, 1.291629431144141e+17, 1.291629431176954e+17, 1.291629431208204e+17, 1.291629431241016e+17, 1.291629431272266e+17, 1.291629431305079e+17, 1.291629431337891e+17, 1.29162943136914e+17, 1.291629431401953e+17, 1.291629431433203e+17, 1.291629431466016e+17, 1.291629431498829e+17, 1.291629431530079e+17, 1.29162943156289e+17, 1.291629431594141e+17, 1.291629431626953e+17, 1.291629431659766e+17, 1.291629431691016e+17, 1.291629431723828e+17, 1.291629431755078e+17, 1.291629431787891e+17, 1.291629431820704e+17, 1.291629431851954e+17, 1.291629431884765e+17, 1.291629431916015e+17, 1.291629431948828e+17, 1.291629431981641e+17, 1.291629432012891e+17, 1.291629432045704e+17, 1.291629432076954e+17, 1.291629432109765e+17, 1.291629432142579e+17, 1.291629432173828e+17, 1.291629432206641e+17, 1.291629432237891e+17, 1.291629432270703e+17, 1.291629432303516e+17, 1.291629432334766e+17, 1.291629432367579e+17, 1.291629432398829e+17, 1.29162943243164e+17, 1.291629432464454e+17, 1.291629432495703e+17, 1.291629432528516e+17, 1.291629432559766e+17, 1.291629432592579e+17, 1.29162943262539e+17, 1.291629432656641e+17, 1.291629432689454e+17, 1.291629432722266e+17, 1.291629432753516e+17, 1.29162943278633e+17, 1.291629432817578e+17, 1.291629432850391e+17, 1.291629432881641e+17, 1.291629432914454e+17, 1.291629432947265e+17, 1.291629432978515e+17, 1.291629433011329e+17, 1.291629433042578e+17, 1.291629433075391e+17, 1.291629433108204e+17, 1.291629433139453e+17, 1.291629433172265e+17, 1.291629433203516e+17, 1.291629433236329e+17, 1.29162943326914e+17, 1.29162943330039e+17, 1.291629433333204e+17, 1.291629433364453e+17, 1.291629433397266e+17, 1.291629433430079e+17, 1.291629433461329e+17, 1.29162943349414e+17, 1.29162943352539e+17, 1.291629433558204e+17, 1.291629433591016e+17, 1.291629433622266e+17, 1.291629433655078e+17, 1.291629433686328e+17, 1.291629433719141e+17, 1.291629433751954e+17, 1.291629433783204e+17, 1.291629433816015e+17, 1.291629433848829e+17, 1.291629433880079e+17, 1.291629433912891e+17, 1.291629433944141e+17, 1.291629433976954e+17, 1.291629434009766e+17, 1.291629434041015e+17, 1.291629434073829e+17, 1.291629434105079e+17, 1.291629434137891e+17, 1.291629434170703e+17, 1.291629434201955e+17, 1.291629434234766e+17, 1.291629434266016e+17, 1.291629434298829e+17, 1.291629434331642e+17, 1.29162943436289e+17, 1.291629434395704e+17, 1.291629434428516e+17, 1.291629434459766e+17, 1.291629434492579e+17, 1.291629434523828e+17, 1.291629434556641e+17, 1.291629434589454e+17, 1.291629434620704e+17, 1.291629434653516e+17, 1.291629434684765e+17, 1.291629434717578e+17, 1.291629434750391e+17, 1.291629434781641e+17, 1.291629434814454e+17, 1.291629434847265e+17, 1.291629434878516e+17, 1.291629434911328e+17, 1.291629434942579e+17, 1.291629434975391e+17, 1.291629435008204e+17, 1.291629435039453e+17, 1.291629435072266e+17, 1.291629435103516e+17, 1.291629435136329e+17, 1.29162943516914e+17, 1.29162943520039e+17, 1.291629435233203e+17, 1.291629435266016e+17, 1.291629435297266e+17, 1.291629435330079e+17, 1.291629435361329e+17, 1.291629435394141e+17, 1.291629435426953e+17, 1.291629435458204e+17, 1.291629435491016e+17, 1.291629435522266e+17, 1.291629435555078e+17, 1.291629435586328e+17, 1.291629435619141e+17, 1.291629435651953e+17, 1.291629435683204e+17, 1.291629435716015e+17, 1.291629435748828e+17, 1.291629435780078e+17, 1.291629435812891e+17, 1.291629435844141e+17, 1.291629435876954e+17, 1.291629435908204e+17, 1.291629435941016e+17, 1.291629435973828e+17, 1.291629436005079e+17, 1.291629436037891e+17, 1.29162943606914e+17, 1.291629436101953e+17, 1.291629436134766e+17, 1.291629436166016e+17, 1.291629436198829e+17, 1.291629436231642e+17, 1.29162943626289e+17, 1.291629436295703e+17, 1.291629436326954e+17, 1.291629436359766e+17, 1.291629436391016e+17, 1.291629436423828e+17, 1.291629436456641e+17, 1.291629436487891e+17, 1.291629436520703e+17, 1.291629436551954e+17, 1.291629436584765e+17, 1.291629436617578e+17, 1.291629436648828e+17, 1.291629436681641e+17, 1.291629436712891e+17, 1.291629436745704e+17, 1.291629436778516e+17, 1.291629436809766e+17, 1.291629436842578e+17, 1.291629436873829e+17, 1.291629436906641e+17, 1.291629436939453e+17, 1.291629436970703e+17, 1.291629437003516e+17, 1.291629437034766e+17, 1.291629437067579e+17, 1.291629437100392e+17, 1.29162943713164e+17, 1.291629437164453e+17, 1.291629437197266e+17, 1.291629437228516e+17, 1.291629437261327e+17, 1.291629437292579e+17, 1.291629437325391e+17, 1.291629437358203e+17, 1.291629437389453e+17, 1.291629437422267e+17, 1.291629437455078e+17, 1.291629437486328e+17, 1.291629437519141e+17, 1.291629437550391e+17, 1.291629437583203e+17, 1.291629437614454e+17, 1.291629437647267e+17, 1.291629437680078e+17, 1.291629437711328e+17, 1.291629437744141e+17, 1.291629437776954e+17, 1.291629437808204e+17, 1.291629437841016e+17, 1.291629437872266e+17, 1.291629437905078e+17, 1.291629437937892e+17, 1.291629437969142e+17, 1.291629438001953e+17, 1.291629438033203e+17, 1.291629438066016e+17, 1.291629438098829e+17, 1.291629438130077e+17, 1.291629438162892e+17, 1.291629438194141e+17, 1.291629438226953e+17, 1.291629438258203e+17, 1.291629438291017e+17, 1.291629438323828e+17, 1.291629438355078e+17, 1.291629438387891e+17, 1.291629438420704e+17, 1.291629438451953e+17, 1.291629438484767e+17, 1.291629438516017e+17, 1.291629438548828e+17, 1.291629438581641e+17, 1.291629438612891e+17, 1.291629438645704e+17, 1.291629438676952e+17, 1.291629438709766e+17, 1.291629438742578e+17, 1.291629438773828e+17, 1.291629438806641e+17, 1.291629438837892e+17, 1.291629438870703e+17, 1.291629438903516e+17, 1.291629438934766e+17, 1.291629438967579e+17, 1.291629438998828e+17, 1.291629439031642e+17, 1.291629439064453e+17, 1.291629439095703e+17, 1.291629439128516e+17, 1.291629439159766e+17, 1.291629439192579e+17, 1.291629439225391e+17, 1.291629439256641e+17, 1.291629439289453e+17, 1.291629439320703e+17, 1.291629439353517e+17, 1.291629439386328e+17, 1.291629439417578e+17, 1.291629439450391e+17, 1.291629439483204e+17, 1.291629439514454e+17, 1.291629439547267e+17, 1.291629439578516e+17, 1.291629439611328e+17, 1.291629439644141e+17, 1.291629439675391e+17, 1.291629439708204e+17, 1.291629439739453e+17, 1.291629439772266e+17, 1.291629439805078e+17, 1.291629439836329e+17, 1.291629439869142e+17, 1.291629439901953e+17, 1.291629439933203e+17, 1.291629439966016e+17, 1.291629439997266e+17, 1.291629440030079e+17, 1.291629440062892e+17, 1.291629440094141e+17, 1.291629440126953e+17, 1.291629440158203e+17, 1.291629440191017e+17, 1.291629440223828e+17, 1.291629440255078e+17, 1.291629440287891e+17, 1.291629440319141e+17, 1.291629440351953e+17, 1.291629440384765e+17, 1.291629440416017e+17, 1.291629440448828e+17, 1.291629440480078e+17, 1.291629440512891e+17, 1.291629440545704e+17, 1.291629440576954e+17, 1.291629440609766e+17, 1.291629440641016e+17, 1.291629440673828e+17, 1.291629440706641e+17, 1.291629440737892e+17, 1.291629440770703e+17, 1.291629440801953e+17, 1.291629440834766e+17, 1.291629440867579e+17, 1.291629440898829e+17, 1.291629440931642e+17, 1.291629440962892e+17, 1.291629440995703e+17, 1.291629441028516e+17, 1.291629441059767e+17, 1.291629441092579e+17, 1.291629441123828e+17, 1.291629441156641e+17, 1.291629441189454e+17, 1.291629441220703e+17, 1.291629441253516e+17, 1.291629441286328e+17, 1.291629441317578e+17, 1.291629441350391e+17, 1.291629441381641e+17, 1.291629441414454e+17, 1.291629441447265e+17, 1.291629441478516e+17, 1.291629441511329e+17, 1.291629441542578e+17, 1.291629441575391e+17, 1.291629441608204e+17, 1.291629441639453e+17, 1.291629441672266e+17, 1.291629441703516e+17, 1.291629441736329e+17, 1.29162944176914e+17, 1.291629441800392e+17, 1.291629441833203e+17, 1.291629441864453e+17, 1.291629441897266e+17, 1.291629441928516e+17, 1.291629441961329e+17, 1.29162944199414e+17, 1.291629442025391e+17, 1.291629442058204e+17, 1.291629442089453e+17, 1.291629442122266e+17, 1.291629442155078e+17, 1.291629442186328e+17, 1.291629442219141e+17, 1.291629442250391e+17, 1.291629442283204e+17, 1.291629442316015e+17, 1.291629442347267e+17, 1.291629442380079e+17, 1.291629442411328e+17, 1.291629442444141e+17, 1.291629442476954e+17, 1.291629442508204e+17, 1.291629442541015e+17, 1.291629442572266e+17, 1.291629442605079e+17, 1.291629442636328e+17, 1.29162944266914e+17, 1.291629442701953e+17, 1.291629442733203e+17, 1.291629442766016e+17, 1.291629442798829e+17, 1.291629442830079e+17, 1.29162944286289e+17, 1.291629442894141e+17, 1.291629442926954e+17, 1.291629442959766e+17, 1.291629442991016e+17, 1.291629443023828e+17, 1.291629443055078e+17, 1.291629443087891e+17, 1.291629443120704e+17, 1.291629443151954e+17, 1.291629443184765e+17, 1.291629443216017e+17, 1.291629443248828e+17, 1.291629443281641e+17, 1.291629443312891e+17, 1.291629443345704e+17, 1.291629443376954e+17, 1.291629443409765e+17, 1.291629443442579e+17, 1.291629443473829e+17, 1.291629443506641e+17, 1.291629443537891e+17, 1.291629443570703e+17, 1.291629443603516e+17, 1.291629443634766e+17, 1.291629443667579e+17, 1.291629443698829e+17, 1.29162944373164e+17, 1.291629443764453e+17, 1.291629443795704e+17, 1.291629443828516e+17, 1.291629443859766e+17, 1.291629443892579e+17, 1.291629443923828e+17, 1.291629443956641e+17, 1.291629443989454e+17, 1.291629444020704e+17, 1.291629444053516e+17, 1.291629444086328e+17, 1.291629444117578e+17, 1.291629444150391e+17, 1.291629444181641e+17, 1.291629444214454e+17, 1.291629444247265e+17, 1.291629444278515e+17, 1.291629444311328e+17, 1.291629444342579e+17, 1.291629444375391e+17, 1.291629444408204e+17, 1.291629444439453e+17, 1.291629444472266e+17, 1.291629444503516e+17, 1.291629444536329e+17, 1.29162944456914e+17, 1.29162944460039e+17, 1.291629444633203e+17, 1.291629444666016e+17, 1.291629444697266e+17, 1.291629444730079e+17, 1.291629444761329e+17, 1.29162944479414e+17, 1.291629444826954e+17, 1.291629444858204e+17, 1.291629444891016e+17, 1.291629444922266e+17, 1.291629444955078e+17, 1.291629444987891e+17, 1.291629445019141e+17, 1.291629445051954e+17, 1.291629445083204e+17, 1.291629445116015e+17, 1.291629445148829e+17, 1.291629445180078e+17, 1.291629445212891e+17, 1.291629445244141e+17, 1.291629445276954e+17, 1.291629445309765e+17, 1.291629445341016e+17, 1.291629445373829e+17, 1.291629445405079e+17, 1.291629445437891e+17, 1.291629445470705e+17, 1.291629445501953e+17, 1.291629445534766e+17, 1.291629445566016e+17, 1.291629445598829e+17, 1.29162944563164e+17, 1.29162944566289e+17, 1.291629445695704e+17, 1.291629445728516e+17, 1.291629445759766e+17, 1.291629445792579e+17, 1.291629445823828e+17, 1.29162944585664e+17, 1.291629445889454e+17, 1.291629445920704e+17, 1.291629445953516e+17, 1.291629445984765e+17, 1.29162944601758e+17, 1.291629446050391e+17, 1.291629446081641e+17, 1.291629446114454e+17, 1.291629446145704e+17, 1.291629446178515e+17, 1.291629446211329e+17, 1.291629446242579e+17, 1.291629446275391e+17, 1.291629446306641e+17, 1.291629446339455e+17, 1.291629446372266e+17, 1.291629446403516e+17, 1.291629446436329e+17, 1.291629446469142e+17, 1.29162944650039e+17, 1.291629446533203e+17, 1.291629446564454e+17, 1.291629446597266e+17, 1.291629446630079e+17, 1.291629446661329e+17, 1.291629446694141e+17, 1.29162944672539e+17, 1.291629446758204e+17, 1.291629446791016e+17, 1.291629446822266e+17, 1.291629446855078e+17, 1.29162944688633e+17, 1.291629446919141e+17, 1.291629446951954e+17, 1.291629446983204e+17, 1.291629447016017e+17, 1.291629447047265e+17, 1.291629447080079e+17, 1.291629447111329e+17, 1.291629447144141e+17, 1.291629447176954e+17, 1.291629447208204e+17, 1.291629447241016e+17, 1.291629447273828e+17, 1.291629447305079e+17, 1.291629447337891e+17, 1.29162944736914e+17, 1.291629447401953e+17, 1.291629447434766e+17, 1.291629447466016e+17, 1.291629447498829e+17, 1.29162944753164e+17, 1.291629447562892e+17, 1.291629447595703e+17, 1.291629447626954e+17, 1.291629447659766e+17, 1.291629447692579e+17, 1.291629447723828e+17, 1.291629447756641e+17, 1.291629447787891e+17, 1.291629447820704e+17, 1.291629447853516e+17, 1.291629447884767e+17, 1.291629447917578e+17, 1.291629447948829e+17, 1.291629447981641e+17, 1.291629448014454e+17, 1.291629448045704e+17, 1.291629448078516e+17, 1.291629448109766e+17, 1.291629448142578e+17, 1.291629448175391e+17, 1.291629448206641e+17, 1.291629448239453e+17, 1.291629448270703e+17, 1.291629448303516e+17, 1.291629448336328e+17, 1.291629448367579e+17, 1.29162944840039e+17, 1.291629448431642e+17, 1.291629448464453e+17, 1.291629448497266e+17, 1.291629448528516e+17, 1.291629448561329e+17, 1.291629448592579e+17, 1.291629448625391e+17, 1.291629448658203e+17, 1.291629448689454e+17, 1.291629448722266e+17, 1.291629448753516e+17, 1.291629448786328e+17, 1.291629448819141e+17, 1.291629448850391e+17, 1.291629448883203e+17, 1.291629448914454e+17, 1.291629448947267e+17, 1.291629448980078e+17, 1.291629449011328e+17, 1.291629449044141e+17, 1.291629449075391e+17, 1.291629449108204e+17, 1.291629449141016e+17, 1.291629449172266e+17, 1.291629449205078e+17, 1.291629449236329e+17, 1.29162944926914e+17, 1.291629449301953e+17, 1.291629449333203e+17, 1.291629449366016e+17, 1.291629449397266e+17, 1.291629449430079e+17, 1.291629449462892e+17, 1.291629449494141e+17, 1.291629449526953e+17, 1.291629449558203e+17, 1.291629449591016e+17, 1.291629449623828e+17, 1.291629449655078e+17, 1.291629449687891e+17, 1.291629449719141e+17, 1.291629449751953e+17, 1.291629449784767e+17, 1.291629449816015e+17, 1.291629449848828e+17, 1.291629449881641e+17, 1.291629449912891e+17, 1.291629449945702e+17, 1.291629449976954e+17, 1.291629450009766e+17, 1.291629450042578e+17, 1.291629450073828e+17, 1.291629450106642e+17, 1.291629450137891e+17, 1.291629450170703e+17, 1.291629450201953e+17, 1.291629450234766e+17, 1.291629450267578e+17, 1.291629450298828e+17, 1.291629450331642e+17, 1.291629450362892e+17, 1.291629450395703e+17, 1.291629450428516e+17, 1.291629450459766e+17, 1.291629450492579e+17, 1.291629450523828e+17, 1.291629450556641e+17, 1.291629450589453e+17, 1.291629450620703e+17, 1.291629450653517e+17, 1.291629450684765e+17, 1.291629450717578e+17, 1.291629450748828e+17, 1.291629450781641e+17, 1.291629450814452e+17, 1.291629450847267e+17, 1.291629450878516e+17, 1.291629450911328e+17, 1.291629450944141e+17, 1.291629450975392e+17, 1.291629451008204e+17, 1.291629451039453e+17, 1.291629451072266e+17, 1.291629451105079e+17, 1.291629451136328e+17, 1.291629451169142e+17, 1.291629451200392e+17, 1.291629451233203e+17, 1.291629451264453e+17, 1.291629451297266e+17, 1.291629451330079e+17, 1.291629451361327e+17, 1.291629451394141e+17, 1.291629451426953e+17, 1.291629451458203e+17, 1.291629451491016e+17, 1.291629451522267e+17, 1.291629451555078e+17, 1.291629451587891e+17, 1.291629451619141e+17, 1.291629451651954e+17, 1.291629451683203e+17, 1.291629451716017e+17, 1.291629451748828e+17, 1.291629451780078e+17, 1.291629451812891e+17, 1.291629451844142e+17, 1.291629451876954e+17, 1.291629451909766e+17, 1.291629451941016e+17, 1.291629451973829e+17, 1.291629452005078e+17, 1.291629452037892e+17, 1.291629452070703e+17, 1.291629452101953e+17, 1.291629452134766e+17, 1.291629452166016e+17, 1.291629452198829e+17, 1.291629452231642e+17, 1.291629452262892e+17, 1.291629452295703e+17, 1.291629452326953e+17, 1.291629452359766e+17, 1.291629452392579e+17, 1.291629452423828e+17, 1.291629452456641e+17, 1.291629452487891e+17, 1.291629452520704e+17, 1.291629452553517e+17, 1.291629452584767e+17, 1.291629452617578e+17, 1.291629452648828e+17, 1.291629452681641e+17, 1.291629452714454e+17, 1.291629452745704e+17, 1.291629452778516e+17, 1.291629452809766e+17, 1.291629452842578e+17, 1.291629452875391e+17, 1.291629452906641e+17, 1.291629452939453e+17, 1.291629452970703e+17, 1.291629453003516e+17, 1.291629453036328e+17, 1.291629453067579e+17, 1.291629453100392e+17, 1.291629453131642e+17, 1.291629453164453e+17, 1.291629453197266e+17, 1.291629453228516e+17, 1.291629453261329e+17, 1.291629453294141e+17, 1.291629453325391e+17, 1.291629453358203e+17, 1.291629453389454e+17, 1.291629453422267e+17, 1.291629453455078e+17, 1.291629453486328e+17, 1.291629453519141e+17, 1.291629453550391e+17, 1.291629453583204e+17, 1.291629453614454e+17, 1.291629453647267e+17, 1.291629453680078e+17, 1.291629453711328e+17, 1.291629453744141e+17, 1.291629453776954e+17, 1.291629453808204e+17, 1.291629453841016e+17, 1.291629453872266e+17, 1.291629453905078e+17, 1.291629453936329e+17, 1.291629453969142e+17, 1.291629454001953e+17, 1.291629454033203e+17, 1.291629454066016e+17, 1.291629454098829e+17, 1.291629454130079e+17, 1.29162945416289e+17, 1.291629454194141e+17, 1.291629454226953e+17, 1.291629454258203e+17, 1.291629454291016e+17, 1.291629454323828e+17, 1.291629454355078e+17, 1.291629454387891e+17, 1.291629454419141e+17, 1.291629454451954e+17, 1.291629454484765e+17, 1.291629454516017e+17, 1.291629454548828e+17, 1.291629454580078e+17, 1.291629454612891e+17, 1.291629454645704e+17, 1.291629454676954e+17, 1.291629454709766e+17, 1.291629454741016e+17, 1.291629454773828e+17, 1.291629454806641e+17, 1.291629454837892e+17, 1.291629454870703e+17, 1.291629454903515e+17, 1.291629454934766e+17, 1.291629454967579e+17, 1.291629454998829e+17, 1.29162945503164e+17, 1.291629455064454e+17, 1.291629455095703e+17, 1.291629455128516e+17, 1.291629455159766e+17, 1.291629455192579e+17, 1.29162945522539e+17, 1.291629455256641e+17, 1.291629455289454e+17, 1.291629455320703e+17, 1.291629455353516e+17, 1.291629455386328e+17, 1.291629455417578e+17, 1.291629455450391e+17, 1.291629455481641e+17, 1.291629455514454e+17, 1.291629455547265e+17, 1.291629455578516e+17, 1.291629455611329e+17, 1.291629455644141e+17, 1.291629455675391e+17, 1.291629455708204e+17, 1.291629455739453e+17, 1.291629455772265e+17, 1.291629455805079e+17, 1.291629455836329e+17, 1.29162945586914e+17, 1.29162945590039e+17, 1.291629455933203e+17, 1.291629455964453e+17, 1.291629455997266e+17, 1.291629456030079e+17, 1.291629456061329e+17, 1.29162945609414e+17, 1.291629456126954e+17, 1.291629456158204e+17, 1.291629456191016e+17, 1.291629456222266e+17, 1.291629456255078e+17, 1.291629456286328e+17, 1.291629456319141e+17, 1.291629456351954e+17, 1.291629456383204e+17, 1.291629456416015e+17, 1.291629456448828e+17, 1.291629456480079e+17, 1.291629456512891e+17, 1.291629456544141e+17, 1.291629456576954e+17, 1.291629456609766e+17, 1.291629456641015e+17, 1.291629456673829e+17, 1.291629456705079e+17, 1.291629456737891e+17, 1.291629456770703e+17, 1.291629456801953e+17, 1.291629456834766e+17, 1.291629456866016e+17, 1.291629456898829e+17, 1.29162945693164e+17, 1.29162945696289e+17, 1.291629456995703e+17, 1.291629457026954e+17, 1.291629457059766e+17, 1.291629457092579e+17, 1.291629457123828e+17, 1.291629457156641e+17, 1.291629457189454e+17, 1.291629457220704e+17, 1.291629457253516e+17, 1.291629457284765e+17, 1.291629457317578e+17, 1.291629457348828e+17, 1.291629457381641e+17, 1.291629457414454e+17, 1.291629457445704e+17, 1.291629457478516e+17, 1.291629457509765e+17, 1.291629457542579e+17, 1.291629457575391e+17, 1.291629457606641e+17, 1.291629457639453e+17, 1.291629457672266e+17, 1.291629457703516e+17, 1.291629457736329e+17, 1.291629457767579e+17, 1.29162945780039e+17, 1.291629457833204e+17, 1.291629457864453e+17, 1.291629457897266e+17, 1.291629457930079e+17, 1.291629457961329e+17, 1.29162945799414e+17, 1.291629458025391e+17, 1.291629458058204e+17, 1.291629458089454e+17, 1.291629458122266e+17, 1.291629458155078e+17, 1.291629458186328e+17, 1.291629458219141e+17, 1.291629458251954e+17, 1.291629458283204e+17, 1.291629458316015e+17, 1.291629458347265e+17, 1.291629458380079e+17, 1.291629458412891e+17, 1.291629458444141e+17, 1.291629458476954e+17, 1.291629458508204e+17, 1.291629458541015e+17, 1.291629458573829e+17, 1.291629458605079e+17, 1.291629458637891e+17, 1.29162945866914e+17, 1.291629458701955e+17, 1.291629458734766e+17, 1.291629458766016e+17, 1.291629458798829e+17, 1.291629458831642e+17, 1.29162945886289e+17, 1.291629458895703e+17, 1.291629458926954e+17, 1.291629458959766e+17, 1.291629458992579e+17, 1.291629459023828e+17, 1.291629459056641e+17, 1.291629459087891e+17, 1.291629459120704e+17, 1.291629459153517e+17, 1.291629459184765e+17, 1.291629459217578e+17, 1.291629459248829e+17, 1.291629459281641e+17, 1.291629459314454e+17, 1.291629459345704e+17, 1.291629459378516e+17, 1.291629459409765e+17, 1.291629459442579e+17, 1.291629459473829e+17, 1.291629459506641e+17, 1.291629459539453e+17, 1.291629459570705e+17, 1.291629459603516e+17, 1.291629459636328e+17, 1.291629459667579e+17, 1.291629459700392e+17, 1.29162945973164e+17, 1.291629459764453e+17, 1.291629459797266e+17, 1.291629459828516e+17, 1.291629459861329e+17, 1.291629459892579e+17, 1.291629459925391e+17, 1.291629459958203e+17, 1.291629459989454e+17, 1.291629460022266e+17, 1.291629460055078e+17, 1.291629460086328e+17, 1.291629460119141e+17, 1.291629460150391e+17, 1.291629460183204e+17, 1.291629460214454e+17, 1.291629460247267e+17, 1.291629460280078e+17, 1.291629460311329e+17, 1.291629460344141e+17, 1.291629460376954e+17, 1.291629460408204e+17, 1.291629460441016e+17, 1.291629460472266e+17, 1.291629460505078e+17, 1.291629460537891e+17, 1.291629460569142e+17, 1.291629460601953e+17, 1.291629460633203e+17, 1.291629460666016e+17, 1.291629460698829e+17, 1.291629460730079e+17, 1.291629460762892e+17, 1.291629460794141e+17, 1.291629460826953e+17, 1.291629460859766e+17, 1.291629460891016e+17, 1.291629460923828e+17, 1.291629460955078e+17, 1.291629460987891e+17, 1.291629461020703e+17, 1.291629461051954e+17, 1.291629461084765e+17, 1.291629461116017e+17, 1.291629461148828e+17, 1.291629461181641e+17, 1.291629461212891e+17, 1.291629461245704e+17, 1.291629461276954e+17, 1.291629461309766e+17, 1.291629461342578e+17, 1.291629461373828e+17, 1.291629461406641e+17, 1.291629461437891e+17, 1.291629461470703e+17, 1.291629461503516e+17, 1.291629461534766e+17, 1.291629461567578e+17, 1.291629461598829e+17, 1.291629461631642e+17, 1.291629461664453e+17, 1.291629461695703e+17, 1.291629461728516e+17, 1.291629461759766e+17, 1.291629461792579e+17, 1.291629461823828e+17, 1.291629461856641e+17, 1.291629461889453e+17, 1.291629461920703e+17, 1.291629461953516e+17, 1.291629461986328e+17, 1.291629462017578e+17, 1.291629462050391e+17, 1.291629462081641e+17, 1.291629462114454e+17, 1.291629462147267e+17, 1.291629462178516e+17, 1.291629462211328e+17, 1.291629462242578e+17, 1.291629462275391e+17, 1.291629462308204e+17, 1.291629462339453e+17, 1.291629462372266e+17, 1.291629462403516e+17, 1.291629462436328e+17, 1.291629462469142e+17, 1.29162946250039e+17, 1.291629462533203e+17, 1.291629462566016e+17, 1.291629462597266e+17, 1.291629462630077e+17, 1.291629462661329e+17, 1.291629462694141e+17, 1.291629462726953e+17, 1.291629462758203e+17, 1.291629462791017e+17, 1.291629462822266e+17, 1.291629462855078e+17, 1.291629462887891e+17, 1.291629462919141e+17, 1.291629462951953e+17, 1.291629462983204e+17, 1.291629463016017e+17, 1.291629463048828e+17, 1.291629463080078e+17, 1.291629463112892e+17, 1.291629463144141e+17, 1.291629463176954e+17, 1.291629463209766e+17, 1.291629463241016e+17, 1.291629463273828e+17, 1.291629463305078e+17, 1.291629463337892e+17, 1.291629463370703e+17, 1.291629463401953e+17, 1.291629463434766e+17, 1.291629463466016e+17, 1.291629463498828e+17, 1.291629463531642e+17, 1.291629463562892e+17, 1.291629463595703e+17, 1.291629463626953e+17, 1.291629463659767e+17, 1.291629463692579e+17, 1.291629463723828e+17, 1.291629463756641e+17, 1.291629463789454e+17, 1.291629463820703e+17, 1.291629463853517e+17, 1.291629463884767e+17, 1.291629463917578e+17, 1.291629463948828e+17, 1.291629463981641e+17, 1.291629464014454e+17, 1.291629464045702e+17, 1.291629464078516e+17, 1.291629464109766e+17, 1.291629464142578e+17, 1.291629464175392e+17, 1.291629464206642e+17, 1.291629464239453e+17, 1.291629464270703e+17, 1.291629464303516e+17, 1.291629464336329e+17, 1.291629464367578e+17, 1.291629464400392e+17, 1.291629464431642e+17, 1.291629464464453e+17, 1.291629464497266e+17, 1.291629464528517e+17, 1.291629464561329e+17, 1.291629464594141e+17, 1.291629464625391e+17, 1.291629464658204e+17, 1.291629464689453e+17, 1.291629464722267e+17, 1.291629464755078e+17, 1.291629464786328e+17, 1.291629464819141e+17, 1.291629464850391e+17, 1.291629464883204e+17, 1.291629464914452e+17, 1.291629464947267e+17, 1.291629464980078e+17, 1.291629465011328e+17, 1.291629465044141e+17, 1.291629465076954e+17, 1.291629465108204e+17, 1.291629465141016e+17, 1.291629465172266e+17, 1.291629465205079e+17, 1.291629465237891e+17, 1.291629465269142e+17, 1.291629465301953e+17, 1.291629465333203e+17, 1.291629465366016e+17, 1.291629465398829e+17, 1.291629465430079e+17, 1.291629465462892e+17, 1.291629465494141e+17, 1.291629465526953e+17, 1.291629465559766e+17, 1.291629465591017e+17, 1.291629465623828e+17, 1.291629465655078e+17, 1.291629465687891e+17, 1.291629465720704e+17, 1.291629465751954e+17, 1.291629465784765e+17, 1.291629465816017e+17, 1.291629465848828e+17, 1.291629465881641e+17, 1.291629465912891e+17, 1.291629465945704e+17, 1.291629465978515e+17, 1.291629466009766e+17, 1.291629466042578e+17, 1.291629466073829e+17, 1.291629466106641e+17, 1.291629466139453e+17, 1.291629466170703e+17, 1.291629466203516e+17, 1.291629466234766e+17, 1.291629466267579e+17, 1.29162946630039e+17, 1.291629466331642e+17, 1.291629466364453e+17, 1.291629466395703e+17, 1.291629466428516e+17, 1.291629466461329e+17, 1.291629466492579e+17, 1.29162946652539e+17, 1.291629466556641e+17, 1.291629466589453e+17, 1.291629466620704e+17, 1.291629466653516e+17, 1.291629466686328e+17, 1.291629466717578e+17, 1.291629466750391e+17, 1.291629466783204e+17, 1.291629466814454e+17, 1.291629466847265e+17, 1.291629466878516e+17, 1.291629466911328e+17, 1.291629466944141e+17, 1.291629466975391e+17, 1.291629467008204e+17, 1.291629467039453e+17, 1.291629467072266e+17, 1.291629467105079e+17, 1.291629467136329e+17, 1.29162946716914e+17, 1.291629467201955e+17, 1.291629467233203e+17, 1.291629467266016e+17, 1.291629467297266e+17, 1.291629467330079e+17, 1.291629467361329e+17, 1.29162946739414e+17, 1.291629467426954e+17, 1.291629467458203e+17, 1.291629467491016e+17, 1.291629467522266e+17, 1.291629467555078e+17, 1.29162946758789e+17, 1.291629467619141e+17, 1.291629467651954e+17, 1.291629467684765e+17, 1.291629467716015e+17, 1.291629467748829e+17, 1.291629467780078e+17, 1.291629467812891e+17, 1.291629467844141e+17, 1.291629467876954e+17, 1.291629467909765e+17, 1.291629467941016e+17, 1.291629467973829e+17, 1.291629468006641e+17, 1.291629468037891e+17, 1.291629468070703e+17, 1.291629468101953e+17, 1.291629468134765e+17, 1.291629468167579e+17, 1.291629468198829e+17, 1.29162946823164e+17, 1.29162946826289e+17, 1.291629468295704e+17, 1.291629468328516e+17, 1.291629468359766e+17, 1.291629468392579e+17, 1.291629468423828e+17, 1.29162946845664e+17, 1.291629468489454e+17, 1.291629468520704e+17, 1.291629468553516e+17, 1.291629468584765e+17, 1.29162946861758e+17, 1.291629468650391e+17, 1.291629468681641e+17, 1.291629468714454e+17, 1.291629468745704e+17, 1.291629468778515e+17, 1.291629468811329e+17, 1.291629468842579e+17, 1.291629468875391e+17, 1.291629468906641e+17, 1.291629468939453e+17, 1.291629468972266e+17, 1.291629469003515e+17, 1.291629469036329e+17, 1.291629469067579e+17, 1.29162946910039e+17, 1.291629469133203e+17, 1.291629469164454e+17, 1.291629469197266e+17, 1.291629469228516e+17, 1.291629469261329e+17, 1.291629469294141e+17, 1.29162946932539e+17, 1.291629469358204e+17, 1.291629469389454e+17, 1.291629469422266e+17, 1.291629469455078e+17, 1.291629469486328e+17, 1.291629469519141e+17, 1.29162946955039e+17, 1.291629469583204e+17, 1.291629469616015e+17, 1.291629469647265e+17, 1.291629469680078e+17, 1.291629469711329e+17, 1.291629469744141e+17, 1.291629469776954e+17, 1.291629469808204e+17, 1.291629469841016e+17, 1.291629469872265e+17, 1.291629469905079e+17, 1.291629469937891e+17, 1.29162946996914e+17, 1.291629470001953e+17, 1.291629470033204e+17, 1.291629470066016e+17, 1.291629470098829e+17, 1.291629470130079e+17, 1.291629470162892e+17, 1.29162947019414e+17, 1.291629470226954e+17, 1.291629470259766e+17, 1.291629470291016e+17, 1.291629470323828e+17, 1.291629470355078e+17, 1.291629470387891e+17, 1.291629470420704e+17, 1.291629470451954e+17, 1.291629470484765e+17, 1.291629470516015e+17, 1.291629470548828e+17, 1.291629470581641e+17, 1.291629470612891e+17, 1.291629470645704e+17, 1.291629470676954e+17, 1.291629470709766e+17, 1.291629470742579e+17, 1.291629470773829e+17, 1.291629470806641e+17, 1.291629470839453e+17, 1.291629470870703e+17, 1.291629470903516e+17, 1.291629470934766e+17, 1.291629470967579e+17, 1.291629470998829e+17, 1.29162947103164e+17, 1.291629471064454e+17, 1.291629471095704e+17, 1.291629471128516e+17, 1.291629471159766e+17, 1.291629471192579e+17, 1.291629471225391e+17, 1.291629471256641e+17, 1.291629471289454e+17, 1.291629471322266e+17, 1.291629471353516e+17, 1.291629471386328e+17, 1.291629471419141e+17, 1.291629471450391e+17, 1.291629471483204e+17, 1.291629471514454e+17, 1.291629471547265e+17, 1.291629471580078e+17, 1.291629471611329e+17, 1.291629471644141e+17, 1.291629471676954e+17, 1.291629471708204e+17, 1.291629471741016e+17, 1.291629471772266e+17, 1.291629471805079e+17, 1.291629471837892e+17, 1.29162947186914e+17, 1.291629471901953e+17, 1.291629471933204e+17, 1.291629471966016e+17, 1.291629471998828e+17, 1.291629472030079e+17, 1.291629472062892e+17, 1.29162947209414e+17, 1.291629472126953e+17, 1.291629472159766e+17, 1.291629472191016e+17, 1.291629472223828e+17, 1.291629472255078e+17, 1.291629472287891e+17, 1.291629472320703e+17, 1.291629472351954e+17, 1.291629472384767e+17, 1.291629472416015e+17, 1.291629472448828e+17, 1.291629472481641e+17, 1.291629472512891e+17, 1.291629472545704e+17, 1.291629472576954e+17, 1.291629472609766e+17, 1.291629472642578e+17, 1.291629472673829e+17, 1.291629472706642e+17, 1.291629472737891e+17, 1.291629472770703e+17, 1.291629472803516e+17, 1.291629472834766e+17, 1.291629472867578e+17, 1.291629472898829e+17, 1.291629472931642e+17, 1.291629472964453e+17, 1.291629472995703e+17, 1.291629473028516e+17, 1.291629473059766e+17, 1.291629473092579e+17, 1.291629473125391e+17, 1.291629473156641e+17, 1.291629473189453e+17, 1.291629473220704e+17, 1.291629473253517e+17, 1.291629473286328e+17, 1.291629473317578e+17, 1.291629473350391e+17, 1.291629473381641e+17, 1.291629473414452e+17, 1.291629473445704e+17, 1.291629473478516e+17, 1.291629473511328e+17, 1.291629473542578e+17, 1.291629473575391e+17, 1.291629473608204e+17, 1.291629473639453e+17, 1.291629473672266e+17, 1.291629473703516e+17, 1.291629473736328e+17, 1.29162947376914e+17, 1.291629473800392e+17, 1.291629473833203e+17, 1.291629473864453e+17, 1.291629473897266e+17, 1.291629473930079e+17, 1.291629473961329e+17, 1.291629473994141e+17, 1.291629474026953e+17, 1.291629474058203e+17, 1.291629474091016e+17, 1.291629474122267e+17, 1.291629474155078e+17, 1.291629474186328e+17, 1.291629474219141e+17, 1.291629474251954e+17, 1.291629474283203e+17, 1.291629474316017e+17, 1.291629474347267e+17, 1.291629474380078e+17, 1.291629474412891e+17, 1.291629474444141e+17, 1.291629474476954e+17, 1.291629474509766e+17, 1.291629474541016e+17, 1.291629474573828e+17, 1.291629474605078e+17, 1.291629474637891e+17, 1.291629474670703e+17, 1.291629474701953e+17, 1.291629474734766e+17, 1.291629474766016e+17, 1.291629474798829e+17, 1.291629474831642e+17, 1.291629474862892e+17, 1.291629474895703e+17, 1.291629474928517e+17, 1.291629474959766e+17, 1.291629474992579e+17, 1.291629475023828e+17, 1.291629475056641e+17, 1.291629475089453e+17, 1.291629475120703e+17, 1.291629475153517e+17, 1.291629475184765e+17, 1.291629475217578e+17, 1.291629475248828e+17, 1.291629475281641e+17, 1.291629475314454e+17, 1.291629475345704e+17, 1.291629475378516e+17, 1.291629475411328e+17, 1.291629475442578e+17, 1.291629475475392e+17, 1.291629475508204e+17, 1.291629475539453e+17, 1.291629475572266e+17, 1.291629475603516e+17, 1.291629475636328e+17, 1.291629475669142e+17, 1.291629475700392e+17, 1.291629475733203e+17, 1.291629475766016e+17, 1.291629475797267e+17, 1.291629475830079e+17, 1.291629475861329e+17, 1.291629475894141e+17, 1.291629475926954e+17, 1.291629475958203e+17, 1.291629475991016e+17, 1.291629476023828e+17, 1.291629476055078e+17, 1.291629476087891e+17, 1.291629476119141e+17, 1.291629476151954e+17, 1.291629476184765e+17, 1.291629476216017e+17, 1.291629476248828e+17, 1.291629476280078e+17, 1.291629476312891e+17, 1.291629476345704e+17, 1.291629476376954e+17, 1.291629476409766e+17, 1.291629476441016e+17, 1.291629476473829e+17, 1.291629476506641e+17, 1.291629476537892e+17, 1.291629476570703e+17, 1.291629476601953e+17, 1.291629476634766e+17, 1.291629476667579e+17, 1.291629476698829e+17, 1.29162947673164e+17, 1.291629476762892e+17, 1.291629476795703e+17, 1.291629476828516e+17, 1.291629476859766e+17, 1.291629476892579e+17, 1.291629476923828e+17, 1.291629476956641e+17, 1.291629476989454e+17, 1.291629477020704e+17, 1.291629477053516e+17, 1.291629477084767e+17, 1.291629477117578e+17, 1.291629477150391e+17, 1.291629477181641e+17, 1.291629477214454e+17, 1.291629477245704e+17, 1.291629477278516e+17, 1.291629477311328e+17, 1.291629477342579e+17, 1.291629477375391e+17, 1.291629477406642e+17, 1.291629477439453e+17, 1.291629477472266e+17, 1.291629477503516e+17, 1.291629477536329e+17, 1.291629477567579e+17, 1.29162947760039e+17, 1.291629477633203e+17, 1.291629477664453e+17, 1.291629477697266e+17, 1.291629477730079e+17, 1.291629477761329e+17, 1.29162947779414e+17, 1.291629477825391e+17, 1.291629477858203e+17, 1.291629477891016e+17, 1.291629477922266e+17, 1.291629477955078e+17, 1.291629477986328e+17, 1.291629478019141e+17, 1.291629478051954e+17, 1.291629478083204e+17, 1.291629478116015e+17, 1.291629478147265e+17, 1.291629478180078e+17, 1.291629478212891e+17, 1.291629478244141e+17, 1.291629478276954e+17, 1.291629478309765e+17, 1.291629478341016e+17, 1.291629478373829e+17, 1.291629478405079e+17, 1.291629478437891e+17, 1.291629478470705e+17, 1.291629478501953e+17, 1.291629478534766e+17, 1.291629478566016e+17, 1.291629478598829e+17, 1.291629478630079e+17, 1.29162947866289e+17, 1.291629478695704e+17, 1.291629478726953e+17, 1.291629478759766e+17, 1.291629478792579e+17, 1.291629478823828e+17, 1.29162947885664e+17, 1.291629478887891e+17, 1.291629478920704e+17, 1.291629478953516e+17, 1.291629478984765e+17, 1.29162947901758e+17, 1.291629479048828e+17, 1.291629479081641e+17, 1.291629479114454e+17, 1.291629479145704e+17, 1.291629479178515e+17, 1.291629479209765e+17, 1.291629479242579e+17, 1.291629479275391e+17, 1.291629479306641e+17, 1.291629479339453e+17, 1.291629479370703e+17, 1.291629479403515e+17, 1.291629479436329e+17, 1.291629479467579e+17, 1.29162947950039e+17, 1.29162947953164e+17, 1.291629479564454e+17, 1.291629479597266e+17, 1.291629479628516e+17, 1.291629479661329e+17, 1.291629479692579e+17, 1.29162947972539e+17, 1.291629479758204e+17, 1.291629479789454e+17, 1.291629479822266e+17, 1.291629479853516e+17, 1.29162947988633e+17, 1.291629479919141e+17, 1.291629479950391e+17, 1.291629479983204e+17, 1.291629480014454e+17, 1.291629480047265e+17, 1.291629480080079e+17, 1.291629480111329e+17, 1.291629480144141e+17, 1.291629480176954e+17, 1.291629480208204e+17, 1.291629480241016e+17, 1.291629480273829e+17, 1.291629480305079e+17, 1.291629480337891e+17, 1.29162948036914e+17, 1.291629480401953e+17, 1.291629480434766e+17, 1.291629480466016e+17, 1.291629480498829e+17, 1.291629480530079e+17, 1.291629480562892e+17, 1.29162948059414e+17, 1.291629480626954e+17, 1.291629480659766e+17, 1.291629480691016e+17, 1.291629480723828e+17, 1.291629480755078e+17, 1.291629480787891e+17, 1.291629480820704e+17, 1.291629480851954e+17, 1.291629480884765e+17, 1.291629480916015e+17, 1.291629480948829e+17, 1.291629480981641e+17, 1.291629481012891e+17, 1.291629481045704e+17, 1.291629481076954e+17, 1.291629481109766e+17, 1.291629481142579e+17, 1.291629481173829e+17, 1.291629481206641e+17, 1.291629481237891e+17, 1.291629481270703e+17, 1.291629481303516e+17, 1.291629481334766e+17, 1.291629481367579e+17, 1.291629481398829e+17, 1.291629481431642e+17, 1.291629481464453e+17, 1.291629481495704e+17, 1.291629481528516e+17, 1.291629481559766e+17, 1.291629481592579e+17, 1.291629481623828e+17, 1.291629481656641e+17, 1.291629481689454e+17, 1.291629481722266e+17, 1.291629481753516e+17, 1.291629481786328e+17, 1.291629481817578e+17, 1.291629481850391e+17, 1.291629481883204e+17, 1.291629481914454e+17, 1.291629481947265e+17, 1.291629481980078e+17, 1.291629482011328e+17, 1.291629482044141e+17, 1.291629482075391e+17, 1.291629482108204e+17, 1.291629482139453e+17, 1.291629482172266e+17, 1.291629482205078e+17, 1.291629482236329e+17, 1.29162948226914e+17, 1.29162948230039e+17, 1.291629482333203e+17, 1.291629482366016e+17, 1.291629482397266e+17, 1.291629482430079e+17, 1.291629482461329e+17, 1.291629482494141e+17, 1.291629482526953e+17, 1.291629482558204e+17, 1.291629482591016e+17, 1.291629482622266e+17, 1.291629482655078e+17, 1.291629482687891e+17, 1.291629482719141e+17, 1.291629482751953e+17, 1.291629482783204e+17, 1.291629482816015e+17, 1.291629482848828e+17, 1.291629482880078e+17, 1.291629482912891e+17, 1.291629482944141e+17, 1.291629482976954e+17, 1.291629483009766e+17, 1.291629483041016e+17, 1.291629483073828e+17, 1.291629483106642e+17, 1.291629483137891e+17, 1.291629483170703e+17, 1.291629483201953e+17, 1.291629483234766e+17, 1.291629483266016e+17, 1.291629483298829e+17, 1.291629483331642e+17, 1.29162948336289e+17, 1.291629483395703e+17, 1.291629483426954e+17, 1.291629483459766e+17, 1.291629483492577e+17, 1.291629483523828e+17, 1.291629483556641e+17, 1.291629483587891e+17, 1.291629483620703e+17, 1.291629483653517e+17, 1.291629483684765e+17, 1.291629483717578e+17, 1.291629483748828e+17, 1.291629483781641e+17, 1.291629483814452e+17, 1.291629483845704e+17, 1.291629483878516e+17, 1.291629483909766e+17, 1.291629483942578e+17, 1.291629483975392e+17, 1.291629484006641e+17, 1.291629484039453e+17, 1.291629484070703e+17, 1.291629484103516e+17, 1.291629484136328e+17, 1.291629484167579e+17, 1.291629484200392e+17, 1.29162948423164e+17, 1.291629484264453e+17, 1.291629484297266e+17, 1.291629484328516e+17, 1.291629484361327e+17, 1.291629484392579e+17, 1.291629484425391e+17, 1.291629484458203e+17, 1.291629484489453e+17, 1.291629484522267e+17, 1.291629484553516e+17, 1.291629484586328e+17, 1.291629484619141e+17, 1.291629484650391e+17, 1.291629484683203e+17, 1.291629484716017e+17, 1.291629484747267e+17, 1.291629484780078e+17, 1.291629484811328e+17, 1.291629484844141e+17, 1.291629484876954e+17, 1.291629484908204e+17, 1.291629484941016e+17, 1.291629484972266e+17, 1.291629485005078e+17, 1.291629485037892e+17, 1.291629485069142e+17, 1.291629485101953e+17, 1.291629485134766e+17, 1.291629485166016e+17, 1.291629485198829e+17, 1.291629485231642e+17, 1.291629485262892e+17, 1.291629485295703e+17, 1.291629485326953e+17, 1.291629485359766e+17, 1.291629485392579e+17, 1.291629485423828e+17, 1.291629485456641e+17, 1.291629485487891e+17, 1.291629485520704e+17, 1.291629485551953e+17, 1.291629485584767e+17, 1.291629485617578e+17, 1.291629485648828e+17, 1.291629485681641e+17, 1.291629485714454e+17, 1.291629485745704e+17, 1.291629485778516e+17, 1.291629485809766e+17, 1.291629485842578e+17, 1.291629485875392e+17, 1.291629485906641e+17, 1.291629485939453e+17, 1.291629485970703e+17, 1.291629486003516e+17, 1.291629486036328e+17, 1.291629486067579e+17, 1.291629486100392e+17, 1.291629486131642e+17, 1.291629486164453e+17, 1.291629486197266e+17, 1.291629486228516e+17, 1.291629486261329e+17, 1.291629486292579e+17, 1.291629486325391e+17, 1.291629486358203e+17, 1.291629486389453e+17, 1.291629486422267e+17, 1.291629486453517e+17, 1.291629486486328e+17, 1.291629486519141e+17, 1.291629486550391e+17, 1.291629486583204e+17, 1.291629486614454e+17, 1.291629486647267e+17, 1.291629486680078e+17, 1.291629486711328e+17, 1.291629486744141e+17, 1.291629486775391e+17, 1.291629486808204e+17, 1.291629486841016e+17, 1.291629486872266e+17, 1.291629486905078e+17, 1.291629486936329e+17, 1.291629486969142e+17, 1.291629487001953e+17, 1.291629487033203e+17, 1.291629487066016e+17, 1.291629487097266e+17, 1.291629487130079e+17, 1.291629487162892e+17, 1.291629487194141e+17, 1.291629487226953e+17, 1.291629487258203e+17, 1.291629487291017e+17, 1.291629487323828e+17, 1.291629487355078e+17, 1.291629487387891e+17, 1.291629487419141e+17, 1.291629487451953e+17, 1.291629487484765e+17, 1.291629487516017e+17, 1.291629487548828e+17, 1.291629487580078e+17, 1.291629487612891e+17, 1.291629487644141e+17, 1.291629487676954e+17, 1.291629487709766e+17, 1.291629487741016e+17, 1.291629487773828e+17, 1.291629487805078e+17, 1.291629487837892e+17, 1.291629487870703e+17, 1.291629487901953e+17, 1.291629487934766e+17, 1.291629487966016e+17, 1.291629487998829e+17, 1.291629488031642e+17, 1.291629488062892e+17, 1.291629488095703e+17, 1.291629488126953e+17, 1.291629488159767e+17, 1.291629488192579e+17, 1.291629488223828e+17, 1.291629488256641e+17, 1.291629488289454e+17, 1.291629488320703e+17, 1.291629488353516e+17, 1.291629488384767e+17, 1.291629488417578e+17, 1.291629488450391e+17, 1.291629488481641e+17, 1.291629488514454e+17, 1.291629488545704e+17, 1.291629488578516e+17, 1.291629488611329e+17, 1.291629488642578e+17, 1.291629488675391e+17, 1.291629488708204e+17, 1.291629488739453e+17, 1.291629488772266e+17, 1.291629488803516e+17, 1.291629488836329e+17, 1.29162948886914e+17, 1.291629488900392e+17, 1.291629488933203e+17, 1.291629488964453e+17, 1.291629488997266e+17, 1.291629489030079e+17, 1.291629489061329e+17, 1.29162948909414e+17, 1.291629489126953e+17, 1.291629489158204e+17, 1.291629489191016e+17, 1.291629489222266e+17, 1.291629489255078e+17, 1.291629489286328e+17, 1.291629489319141e+17, 1.291629489351954e+17, 1.291629489383204e+17, 1.291629489416015e+17, 1.291629489448828e+17, 1.291629489480079e+17, 1.291629489512891e+17, 1.291629489544141e+17, 1.291629489576954e+17, 1.291629489609766e+17, 1.291629489641015e+17, 1.291629489673829e+17, 1.291629489705079e+17, 1.291629489737891e+17, 1.291629489770703e+17, 1.291629489801953e+17, 1.291629489834766e+17, 1.291629489866016e+17, 1.291629489898829e+17, 1.29162948993164e+17, 1.29162948996289e+17, 1.291629489995703e+17, 1.291629490026954e+17, 1.291629490059766e+17, 1.291629490092579e+17, 1.291629490123828e+17, 1.291629490156641e+17, 1.291629490187891e+17, 1.291629490220704e+17, 1.291629490253516e+17, 1.291629490284765e+17, 1.291629490317578e+17, 1.291629490348828e+17, 1.291629490381641e+17, 1.291629490414454e+17, 1.291629490445704e+17, 1.291629490478515e+17, 1.291629490509765e+17, 1.291629490542579e+17, 1.291629490573829e+17, 1.291629490606641e+17, 1.291629490639453e+17, 1.291629490670703e+17, 1.291629490703516e+17, 1.291629490736329e+17, 1.291629490767579e+17, 1.29162949080039e+17, 1.29162949083164e+17, 1.291629490864453e+17, 1.291629490897266e+17, 1.291629490928516e+17, 1.291629490961329e+17, 1.291629490992579e+17, 1.291629491025391e+17, 1.291629491058204e+17, 1.291629491089454e+17, 1.291629491122266e+17, 1.291629491153516e+17, 1.291629491186328e+17, 1.291629491219141e+17, 1.291629491250391e+17, 1.291629491283204e+17, 1.291629491314454e+17, 1.291629491347265e+17, 1.291629491380079e+17, 1.291629491411328e+17, 1.291629491444141e+17, 1.291629491475391e+17, 1.291629491508204e+17, 1.291629491541015e+17, 1.291629491572266e+17, 1.291629491605079e+17, 1.291629491636329e+17, 1.29162949166914e+17, 1.291629491701955e+17, 1.291629491733203e+17, 1.291629491766016e+17, 1.291629491798829e+17, 1.291629491830079e+17, 1.29162949186289e+17, 1.29162949189414e+17, 1.291629491926954e+17, 1.291629491959766e+17, 1.291629491991016e+17, 1.291629492023828e+17, 1.291629492056641e+17, 1.291629492087891e+17, 1.291629492120704e+17, 1.291629492151954e+17, 1.291629492184765e+17, 1.291629492217578e+17, 1.291629492248829e+17, 1.291629492281641e+17, 1.291629492312891e+17, 1.291629492345704e+17, 1.291629492378516e+17, 1.291629492409765e+17, 1.291629492442579e+17, 1.291629492473829e+17, 1.291629492506641e+17, 1.291629492539453e+17, 1.291629492570705e+17, 1.291629492603516e+17, 1.291629492634766e+17, 1.291629492667579e+17, 1.291629492700392e+17, 1.29162949273164e+17, 1.291629492764454e+17, 1.291629492795704e+17, 1.291629492828516e+17, 1.291629492861329e+17, 1.291629492892579e+17, 1.291629492925391e+17, 1.29162949295664e+17, 1.291629492989454e+17, 1.291629493022266e+17, 1.291629493053516e+17, 1.291629493086328e+17, 1.291629493119141e+17, 1.291629493150391e+17, 1.291629493183204e+17, 1.291629493214454e+17, 1.291629493247267e+17, 1.291629493280078e+17, 1.291629493311329e+17, 1.291629493344141e+17, 1.291629493375391e+17, 1.291629493408204e+17, 1.291629493441016e+17, 1.291629493472266e+17, 1.291629493505079e+17, 1.291629493536329e+17, 1.291629493569142e+17, 1.291629493601953e+17, 1.291629493633204e+17, 1.291629493666016e+17, 1.291629493697266e+17, 1.291629493730079e+17, 1.291629493762892e+17, 1.291629493794141e+17, 1.291629493826953e+17, 1.291629493858204e+17, 1.291629493891016e+17, 1.291629493923828e+17, 1.291629493955078e+17, 1.291629493987891e+17, 1.291629494019141e+17, 1.291629494051954e+17, 1.291629494084765e+17, 1.291629494116017e+17, 1.291629494148828e+17, 1.291629494180079e+17, 1.291629494212891e+17, 1.291629494244141e+17, 1.291629494276954e+17, 1.291629494309766e+17, 1.291629494341016e+17, 1.291629494373828e+17, 1.291629494406641e+17, 1.291629494437891e+17, 1.291629494470703e+17, 1.291629494501953e+17, 1.291629494534766e+17, 1.291629494566016e+17, 1.291629494598829e+17, 1.29162949463164e+17, 1.291629494662892e+17, 1.291629494695703e+17, 1.291629494726954e+17, 1.291629494759766e+17, 1.291629494792579e+17, 1.291629494823828e+17, 1.291629494856641e+17, 1.291629494887891e+17, 1.291629494920704e+17, 1.291629494953516e+17, 1.291629494984767e+17, 1.291629495017578e+17, 1.291629495048829e+17, 1.291629495081641e+17, 1.291629495114454e+17, 1.291629495145704e+17, 1.291629495178516e+17, 1.291629495209766e+17, 1.291629495242578e+17, 1.291629495275391e+17, 1.291629495306641e+17, 1.291629495339453e+17, 1.291629495372266e+17, 1.291629495403516e+17, 1.291629495436328e+17, 1.291629495467579e+17, 1.29162949550039e+17, 1.291629495533203e+17, 1.291629495564453e+17, 1.291629495597266e+17, 1.291629495628516e+17, 1.291629495661329e+17, 1.291629495694141e+17, 1.291629495725391e+17, 1.291629495758203e+17, 1.291629495789454e+17, 1.291629495822266e+17, 1.291629495855078e+17, 1.291629495886328e+17, 1.291629495919141e+17, 1.291629495950391e+17, 1.291629495983203e+17, 1.291629496016017e+17, 1.291629496047265e+17, 1.291629496080078e+17, 1.291629496111328e+17, 1.291629496144141e+17, 1.291629496176954e+17, 1.291629496208204e+17, 1.291629496241016e+17, 1.291629496272266e+17, 1.291629496305078e+17, 1.291629496337892e+17, 1.29162949636914e+17, 1.291629496401953e+17, 1.291629496433203e+17, 1.291629496466016e+17, 1.291629496498828e+17, 1.291629496530079e+17, 1.291629496562892e+17, 1.291629496594141e+17, 1.291629496626953e+17, 1.291629496659767e+17, 1.291629496691016e+17, 1.291629496723828e+17, 1.291629496755078e+17, 1.291629496787891e+17, 1.291629496820703e+17, 1.291629496851953e+17, 1.291629496884767e+17, 1.291629496916015e+17, 1.291629496948828e+17, 1.291629496981641e+17, 1.291629497012891e+17, 1.291629497045702e+17, 1.291629497076954e+17, 1.291629497109766e+17, 1.291629497142578e+17, 1.291629497173828e+17, 1.291629497206642e+17, 1.291629497237891e+17, 1.291629497270703e+17, 1.291629497303516e+17, 1.291629497334766e+17, 1.291629497367578e+17, 1.291629497398828e+17, 1.291629497431642e+17, 1.291629497464453e+17, 1.291629497495703e+17, 1.291629497528516e+17, 1.291629497559766e+17, 1.291629497592579e+17, 1.291629497625391e+17, 1.291629497656641e+17, 1.291629497689453e+17, 1.291629497720703e+17, 1.291629497753517e+17, 1.291629497786328e+17, 1.291629497817578e+17, 1.291629497850391e+17, 1.291629497881641e+17, 1.291629497914452e+17, 1.291629497947267e+17, 1.291629497978516e+17, 1.291629498011328e+17, 1.291629498042578e+17, 1.291629498075392e+17, 1.291629498108204e+17, 1.291629498139453e+17, 1.291629498172266e+17, 1.291629498203516e+17, 1.291629498236328e+17, 1.291629498269142e+17, 1.291629498300392e+17, 1.291629498333203e+17, 1.291629498364453e+17, 1.291629498397266e+17, 1.291629498430079e+17, 1.291629498461327e+17, 1.291629498494141e+17, 1.291629498526953e+17, 1.291629498558203e+17, 1.291629498591016e+17, 1.291629498622267e+17, 1.291629498655078e+17, 1.291629498687891e+17, 1.291629498719141e+17, 1.291629498751954e+17, 1.291629498783203e+17, 1.291629498816017e+17, 1.291629498848828e+17, 1.291629498880078e+17, 1.291629498912891e+17, 1.291629498945704e+17, 1.291629498976954e+17, 1.291629499009766e+17, 1.291629499041016e+17, 1.291629499073829e+17, 1.291629499106641e+17, 1.291629499137892e+17, 1.291629499170703e+17, 1.291629499201953e+17, 1.291629499234766e+17, 1.291629499267579e+17, 1.291629499298829e+17, 1.291629499331642e+17, 1.291629499362892e+17, 1.291629499395703e+17, 1.291629499428516e+17, 1.291629499459766e+17, 1.291629499492579e+17, 1.291629499523828e+17, 1.291629499556641e+17, 1.291629499589453e+17, 1.291629499620704e+17, 1.291629499653517e+17, 1.291629499684767e+17, 1.291629499717578e+17, 1.291629499750391e+17, 1.291629499781641e+17, 1.291629499814454e+17, 1.291629499845704e+17, 1.291629499878516e+17, 1.291629499911328e+17, 1.291629499942578e+17, 1.291629499975391e+17, 1.291629500006641e+17, 1.291629500039453e+17, 1.291629500072266e+17, 1.291629500103516e+17, 1.291629500136328e+17, 1.291629500167579e+17, 1.291629500200392e+17, 1.291629500233203e+17, 1.291629500264453e+17, 1.291629500297266e+17, 1.291629500328516e+17, 1.291629500361329e+17, 1.291629500394141e+17, 1.291629500425391e+17, 1.291629500458203e+17, 1.291629500489454e+17, 1.291629500522267e+17, 1.291629500555078e+17, 1.291629500586328e+17, 1.291629500619141e+17, 1.291629500650391e+17, 1.291629500683204e+17, 1.291629500716015e+17, 1.291629500747267e+17, 1.291629500780078e+17, 1.291629500811328e+17, 1.291629500844141e+17, 1.291629500876954e+17, 1.291629500908204e+17, 1.291629500941016e+17, 1.291629500972266e+17, 1.291629501005078e+17, 1.291629501037891e+17, 1.291629501069142e+17, 1.291629501101953e+17, 1.291629501133203e+17, 1.291629501166016e+17, 1.291629501198829e+17, 1.291629501230079e+17, 1.291629501262892e+17, 1.291629501295704e+17, 1.291629501326953e+17, 1.291629501359766e+17, 1.291629501391016e+17, 1.291629501423828e+17, 1.29162950145664e+17, 1.291629501487891e+17, 1.291629501520704e+17, 1.291629501551953e+17, 1.291629501584765e+17, 1.291629501617578e+17, 1.291629501648828e+17, 1.291629501681641e+17, 1.291629501712891e+17, 1.291629501745704e+17, 1.291629501778515e+17, 1.291629501809766e+17, 1.291629501842579e+17, 1.291629501873828e+17, 1.291629501906641e+17, 1.291629501939453e+17, 1.291629501970703e+17, 1.291629502003515e+17, 1.291629502034766e+17, 1.291629502067579e+17, 1.291629502098829e+17, 1.29162950213164e+17, 1.291629502164454e+17, 1.291629502195703e+17, 1.291629502228516e+17, 1.291629502261329e+17, 1.291629502292579e+17, 1.29162950232539e+17, 1.291629502358204e+17, 1.291629502389454e+17, 1.291629502422266e+17, 1.291629502453516e+17, 1.291629502486328e+17, 1.291629502517578e+17, 1.291629502550391e+17, 1.291629502583204e+17, 1.291629502614454e+17, 1.291629502647265e+17, 1.291629502680078e+17, 1.291629502711329e+17, 1.291629502744141e+17, 1.291629502775391e+17, 1.291629502808204e+17, 1.291629502841016e+17, 1.291629502872265e+17, 1.291629502905079e+17, 1.291629502936329e+17, 1.29162950296914e+17, 1.291629503001953e+17, 1.291629503033203e+17, 1.291629503066016e+17, 1.291629503097266e+17, 1.291629503130079e+17, 1.29162950316289e+17, 1.29162950319414e+17, 1.291629503226954e+17, 1.291629503258204e+17, 1.291629503291016e+17, 1.291629503323828e+17, 1.291629503355078e+17, 1.291629503387891e+17, 1.291629503419141e+17, 1.291629503451954e+17, 1.291629503484765e+17, 1.291629503516015e+17, 1.291629503548828e+17, 1.291629503581641e+17, 1.291629503612891e+17, 1.291629503645704e+17, 1.291629503676954e+17, 1.291629503709766e+17, 1.291629503742579e+17, 1.291629503773829e+17, 1.291629503806641e+17, 1.291629503837891e+17, 1.291629503870703e+17, 1.291629503903516e+17, 1.291629503934766e+17, 1.291629503967579e+17, 1.291629503998829e+17, 1.29162950403164e+17, 1.291629504064454e+17, 1.291629504095703e+17, 1.291629504128516e+17, 1.291629504159766e+17, 1.291629504192579e+17, 1.29162950422539e+17, 1.291629504256641e+17, 1.291629504289454e+17, 1.291629504320704e+17, 1.291629504353516e+17, 1.29162950438633e+17, 1.291629504417578e+17, 1.291629504450391e+17, 1.291629504481641e+17, 1.291629504514454e+17, 1.291629504547265e+17, 1.291629504578516e+17, 1.291629504611329e+17, 1.291629504642579e+17, 1.291629504675391e+17, 1.291629504708204e+17, 1.291629504739453e+17, 1.291629504772266e+17, 1.291629504803516e+17, 1.291629504836329e+17, 1.29162950486914e+17, 1.29162950490039e+17, 1.291629504933204e+17, 1.291629504964453e+17, 1.291629504997266e+17, 1.291629505030079e+17, 1.291629505061329e+17, 1.29162950509414e+17, 1.291629505125391e+17, 1.291629505158204e+17, 1.291629505191016e+17, 1.291629505222266e+17, 1.29162950525508e+17, 1.291629505286328e+17, 1.291629505319141e+17, 1.291629505351954e+17, 1.291629505383204e+17, 1.291629505416015e+17, 1.291629505447265e+17, 1.291629505480079e+17, 1.291629505512891e+17, 1.291629505544141e+17, 1.291629505576954e+17, 1.291629505609766e+17, 1.291629505641015e+17, 1.291629505673829e+17, 1.291629505705079e+17, 1.291629505737891e+17, 1.291629505770703e+17, 1.291629505801955e+17, 1.291629505834766e+17, 1.291629505866016e+17, 1.291629505898829e+17, 1.291629505930079e+17, 1.29162950596289e+17, 1.291629505995703e+17, 1.291629506026954e+17, 1.291629506059766e+17, 1.291629506092579e+17, 1.291629506123828e+17, 1.291629506156641e+17, 1.291629506187891e+17, 1.291629506220704e+17, 1.291629506253517e+17, 1.291629506284765e+17, 1.291629506317578e+17, 1.291629506348829e+17, 1.291629506381641e+17, 1.291629506414454e+17, 1.291629506445704e+17, 1.291629506478516e+17, 1.291629506509765e+17, 1.291629506542579e+17, 1.291629506575391e+17, 1.291629506606641e+17, 1.291629506639453e+17, 1.291629506670705e+17, 1.291629506703516e+17, 1.291629506736328e+17, 1.291629506767579e+17, 1.291629506800392e+17, 1.29162950683164e+17, 1.291629506864453e+17, 1.291629506897266e+17, 1.291629506928516e+17, 1.291629506961329e+17, 1.291629506992579e+17, 1.291629507025391e+17, 1.291629507058203e+17, 1.291629507089454e+17, 1.291629507122266e+17, 1.291629507153516e+17, 1.291629507186328e+17, 1.291629507219141e+17, 1.291629507250391e+17, 1.291629507283204e+17, 1.291629507314454e+17, 1.291629507347267e+17, 1.291629507380078e+17, 1.291629507411329e+17, 1.291629507444141e+17, 1.291629507476954e+17, 1.291629507508204e+17, 1.291629507541016e+17, 1.291629507572266e+17, 1.291629507605078e+17, 1.291629507637891e+17, 1.291629507669142e+17, 1.291629507701953e+17, 1.291629507733203e+17, 1.291629507766016e+17, 1.291629507798829e+17, 1.291629507830079e+17, 1.291629507862892e+17, 1.291629507894141e+17, 1.291629507926953e+17, 1.291629507959766e+17, 1.291629507991016e+17, 1.291629508023828e+17, 1.291629508055078e+17, 1.291629508087891e+17, 1.291629508119141e+17, 1.291629508151954e+17, 1.291629508184765e+17, 1.291629508216017e+17, 1.291629508248828e+17, 1.291629508280079e+17, 1.291629508312891e+17, 1.291629508345704e+17, 1.291629508376954e+17, 1.291629508409766e+17, 1.291629508441016e+17, 1.291629508473828e+17, 1.291629508506641e+17, 1.291629508537891e+17, 1.291629508570703e+17, 1.291629508601953e+17, 1.291629508634766e+17, 1.291629508667578e+17, 1.291629508698829e+17, 1.291629508731642e+17, 1.291629508762892e+17, 1.291629508795703e+17, 1.291629508828516e+17, 1.291629508859766e+17, 1.291629508892579e+17, 1.291629508923828e+17, 1.291629508956641e+17, 1.291629508989453e+17, 1.291629509020704e+17, 1.291629509053516e+17, 1.291629509086328e+17, 1.291629509117578e+17, 1.291629509150391e+17, 1.291629509181641e+17, 1.291629509214454e+17, 1.291629509247267e+17, 1.291629509278516e+17, 1.291629509311328e+17, 1.291629509342578e+17, 1.291629509375391e+17, 1.291629509408204e+17, 1.291629509439453e+17, 1.291629509472266e+17, 1.291629509503516e+17, 1.291629509536328e+17, 1.291629509569142e+17, 1.29162950960039e+17, 1.291629509633203e+17, 1.291629509664453e+17, 1.291629509697266e+17, 1.291629509730077e+17, 1.291629509761329e+17, 1.291629509794141e+17, 1.291629509825391e+17, 1.291629509858203e+17, 1.291629509891017e+17, 1.291629509922266e+17, 1.291629509955078e+17, 1.291629509986328e+17, 1.291629510019141e+17, 1.291629510051953e+17, 1.291629510083203e+17, 1.291629510116017e+17, 1.291629510148828e+17, 1.291629510180078e+17, 1.291629510212892e+17, 1.291629510244141e+17, 1.291629510276954e+17, 1.291629510309766e+17, 1.291629510341016e+17, 1.291629510373828e+17, 1.291629510405078e+17, 1.291629510437892e+17, 1.291629510470703e+17, 1.291629510501953e+17, 1.291629510534766e+17, 1.291629510566016e+17, 1.291629510598828e+17, 1.291629510631642e+17, 1.291629510662892e+17, 1.291629510695703e+17, 1.291629510726953e+17, 1.291629510759767e+17, 1.291629510792579e+17, 1.291629510823828e+17, 1.291629510856641e+17, 1.291629510887891e+17, 1.291629510920703e+17, 1.291629510953517e+17, 1.291629510984767e+17, 1.291629511017578e+17, 1.291629511048828e+17, 1.291629511081641e+17, 1.291629511114454e+17, 1.291629511145702e+17, 1.291629511178516e+17, 1.291629511209766e+17, 1.291629511242578e+17, 1.291629511275391e+17, 1.291629511306642e+17, 1.291629511339453e+17, 1.291629511370703e+17, 1.291629511403516e+17, 1.291629511436329e+17, 1.291629511467578e+17, 1.291629511500392e+17, 1.291629511531642e+17, 1.291629511564453e+17, 1.291629511597266e+17, 1.291629511628517e+17, 1.291629511661329e+17, 1.291629511692579e+17, 1.291629511725391e+17, 1.291629511758204e+17, 1.291629511789453e+17, 1.291629511822267e+17, 1.291629511853517e+17, 1.291629511886328e+17, 1.291629511919141e+17, 1.291629511950391e+17, 1.291629511983204e+17, 1.291629512016017e+17, 1.291629512047267e+17, 1.291629512080078e+17, 1.291629512111328e+17, 1.291629512144141e+17, 1.291629512176954e+17, 1.291629512208204e+17, 1.291629512241016e+17, 1.291629512272266e+17, 1.291629512305079e+17, 1.291629512336328e+17, 1.291629512369142e+17, 1.291629512401953e+17, 1.291629512434766e+17, 1.291629512466016e+17, 1.291629512498829e+17, 1.291629512530079e+17, 1.291629512562892e+17, 1.291629512595703e+17, 1.291629512626953e+17, 1.291629512659766e+17, 1.291629512692579e+17, 1.291629512723828e+17, 1.291629512756641e+17, 1.291629512789454e+17, 1.291629512820704e+17, 1.291629512853516e+17, 1.291629512884767e+17, 1.291629512917578e+17, 1.291629512948828e+17, 1.291629512981641e+17, 1.291629513014454e+17, 1.291629513045704e+17, 1.291629513078515e+17, 1.291629513111329e+17, 1.291629513142578e+17, 1.291629513175391e+17, 1.291629513206641e+17, 1.291629513239453e+17, 1.291629513272265e+17, 1.291629513303516e+17, 1.291629513336329e+17, 1.291629513367579e+17, 1.29162951340039e+17, 1.291629513433204e+17, 1.291629513464453e+17, 1.291629513497266e+17, 1.291629513530079e+17, 1.291629513561329e+17, 1.29162951359414e+17, 1.29162951362539e+17, 1.291629513658204e+17, 1.291629513689453e+17, 1.291629513722266e+17, 1.291629513755078e+17, 1.291629513786328e+17, 1.29162951381914e+17, 1.291629513850391e+17, 1.291629513883204e+17, 1.291629513916015e+17, 1.291629513947265e+17, 1.291629513980079e+17, 1.291629514011328e+17, 1.291629514044141e+17, 1.291629514076954e+17, 1.291629514108204e+17, 1.291629514141015e+17, 1.291629514173829e+17, 1.291629514205079e+17, 1.291629514237891e+17, 1.29162951426914e+17, 1.291629514301953e+17, 1.291629514334766e+17, 1.291629514366016e+17, 1.291629514398829e+17, 1.291629514430079e+17, 1.29162951446289e+17, 1.291629514495704e+17, 1.291629514526954e+17, 1.291629514559766e+17, 1.291629514591016e+17, 1.291629514623828e+17, 1.291629514655078e+17, 1.29162951468789e+17, 1.291629514720704e+17, 1.291629514751954e+17, 1.291629514784765e+17, 1.291629514816015e+17, 1.291629514848829e+17, 1.291629514881641e+17, 1.291629514912891e+17, 1.291629514945704e+17, 1.291629514976954e+17, 1.291629515009765e+17, 1.291629515042579e+17, 1.291629515073829e+17, 1.291629515106641e+17, 1.291629515139453e+17, 1.291629515170703e+17, 1.291629515203516e+17, 1.291629515234765e+17, 1.291629515267579e+17, 1.291629515298829e+17, 1.29162951533164e+17, 1.291629515364453e+17, 1.291629515395704e+17, 1.291629515428516e+17, 1.291629515459766e+17, 1.291629515492579e+17, 1.291629515525391e+17, 1.29162951555664e+17, 1.291629515589454e+17, 1.291629515620704e+17, 1.291629515653516e+17, 1.291629515686328e+17, 1.29162951571758e+17, 1.291629515750391e+17, 1.291629515781641e+17, 1.291629515814454e+17, 1.291629515847267e+17, 1.291629515878515e+17, 1.291629515911329e+17, 1.291629515944141e+17, 1.291629515975391e+17, 1.291629516008204e+17, 1.291629516039453e+17, 1.291629516072266e+17, 1.291629516105079e+17, 1.291629516136329e+17, 1.29162951616914e+17, 1.29162951620039e+17, 1.291629516233203e+17, 1.291629516264454e+17, 1.291629516297266e+17, 1.291629516330079e+17, 1.291629516361329e+17, 1.291629516394141e+17, 1.291629516426954e+17, 1.291629516458204e+17, 1.291629516491016e+17, 1.291629516522266e+17, 1.291629516555078e+17, 1.291629516586328e+17, 1.291629516619141e+17, 1.291629516651954e+17, 1.291629516683204e+17, 1.291629516716015e+17, 1.291629516748829e+17, 1.291629516780078e+17, 1.291629516812891e+17, 1.291629516844141e+17, 1.291629516876954e+17, 1.291629516908204e+17, 1.291629516941016e+17, 1.291629516973829e+17, 1.291629517005079e+17, 1.291629517037891e+17, 1.29162951706914e+17, 1.291629517101953e+17, 1.291629517134766e+17, 1.291629517166016e+17, 1.291629517198829e+17, 1.291629517230079e+17, 1.291629517262892e+17, 1.291629517295704e+17, 1.291629517326954e+17, 1.291629517359766e+17, 1.291629517391016e+17, 1.291629517423828e+17, 1.291629517456641e+17, 1.291629517487891e+17, 1.291629517520704e+17, 1.291629517551954e+17, 1.291629517584765e+17, 1.291629517617578e+17, 1.291629517648828e+17, 1.291629517681641e+17, 1.291629517712891e+17, 1.291629517745704e+17, 1.291629517778515e+17, 1.291629517809766e+17, 1.291629517842579e+17, 1.291629517873829e+17, 1.291629517906641e+17, 1.291629517939453e+17, 1.291629517970703e+17, 1.291629518003516e+17, 1.291629518034766e+17, 1.291629518067579e+17, 1.29162951810039e+17, 1.29162951813164e+17, 1.291629518164454e+17, 1.291629518195703e+17, 1.291629518228516e+17, 1.291629518261329e+17, 1.291629518292579e+17, 1.291629518325391e+17, 1.291629518356641e+17, 1.291629518389454e+17, 1.291629518422266e+17, 1.291629518453516e+17, 1.291629518486328e+17, 1.291629518517578e+17, 1.291629518550391e+17, 1.291629518583204e+17, 1.291629518614454e+17, 1.291629518647265e+17, 1.291629518678516e+17, 1.291629518711329e+17, 1.291629518744141e+17, 1.291629518775391e+17, 1.291629518808204e+17, 1.291629518841016e+17, 1.291629518872266e+17, 1.291629518905079e+17, 1.291629518936329e+17, 1.29162951896914e+17, 1.291629519001953e+17, 1.291629519033204e+17, 1.291629519066016e+17, 1.291629519097266e+17, 1.291629519130079e+17, 1.291629519162892e+17, 1.29162951919414e+17, 1.291629519226953e+17, 1.291629519259766e+17, 1.291629519291016e+17, 1.291629519323828e+17, 1.291629519355078e+17, 1.291629519387891e+17, 1.291629519420703e+17, 1.291629519451954e+17, 1.291629519484767e+17, 1.291629519516015e+17, 1.291629519548828e+17, 1.291629519580079e+17, 1.291629519612891e+17, 1.291629519645704e+17, 1.291629519676954e+17, 1.291629519709766e+17, 1.291629519741016e+17, 1.291629519773829e+17, 1.291629519806641e+17, 1.291629519837891e+17, 1.291629519870703e+17, 1.291629519901955e+17, 1.291629519934766e+17, 1.291629519967578e+17, 1.291629519998829e+17, 1.291629520031642e+17, 1.29162952006289e+17, 1.291629520095703e+17, 1.291629520128516e+17, 1.291629520159766e+17, 1.291629520192579e+17, 1.291629520223828e+17, 1.291629520256641e+17, 1.291629520289453e+17, 1.291629520320704e+17, 1.291629520353517e+17, 1.291629520386328e+17, 1.291629520417578e+17, 1.291629520450391e+17, 1.291629520481641e+17, 1.291629520514454e+17, 1.291629520547267e+17, 1.291629520578516e+17, 1.291629520611328e+17, 1.291629520644141e+17, 1.291629520675391e+17, 1.291629520708204e+17, 1.291629520739453e+17, 1.291629520772266e+17, 1.291629520803516e+17, 1.291629520836328e+17, 1.29162952086914e+17, 1.291629520900392e+17, 1.291629520933203e+17, 1.291629520964453e+17, 1.291629520997266e+17, 1.291629521030079e+17, 1.291629521061329e+17, 1.291629521094141e+17, 1.291629521125391e+17, 1.291629521158203e+17, 1.291629521191016e+17, 1.291629521222267e+17, 1.291629521255078e+17, 1.291629521286328e+17, 1.291629521319141e+17, 1.291629521351954e+17, 1.291629521383203e+17, 1.291629521416017e+17, 1.291629521447267e+17, 1.291629521480078e+17, 1.291629521512891e+17, 1.291629521544141e+17, 1.291629521576954e+17, 1.291629521608204e+17, 1.291629521641016e+17, 1.291629521673828e+17, 1.291629521705078e+17, 1.291629521737891e+17, 1.291629521769142e+17, 1.291629521801953e+17, 1.291629521834766e+17, 1.291629521866016e+17, 1.291629521898829e+17, 1.291629521930079e+17, 1.291629521962892e+17, 1.291629521995703e+17, 1.291629522026953e+17, 1.291629522059766e+17, 1.291629522091016e+17, 1.291629522123828e+17, 1.291629522156641e+17, 1.291629522187891e+17, 1.291629522220703e+17, 1.291629522251953e+17, 1.291629522284765e+17, 1.291629522317578e+17, 1.291629522348828e+17, 1.291629522381641e+17, 1.291629522414452e+17, 1.291629522445704e+17, 1.291629522478516e+17, 1.291629522509766e+17, 1.291629522542578e+17, 1.291629522573828e+17, 1.291629522606641e+17, 1.291629522639453e+17, 1.291629522670703e+17, 1.291629522703516e+17, 1.291629522736328e+17, 1.291629522769142e+17, 1.291629522800392e+17, 1.291629522833203e+17, 1.291629522864453e+17, 1.291629522897267e+17, 1.291629522928516e+17, 1.291629522961329e+17, 1.291629522994141e+17, 1.291629523025391e+17, 1.291629523058203e+17, 1.291629523089453e+17, 1.291629523122267e+17, 1.291629523155078e+17, 1.291629523186328e+17, 1.291629523219141e+17, 1.291629523250391e+17, 1.291629523283203e+17, 1.291629523316017e+17, 1.291629523347267e+17, 1.291629523380078e+17, 1.291629523411328e+17, 1.291629523444142e+17, 1.291629523476954e+17, 1.291629523508204e+17, 1.291629523541016e+17, 1.291629523572266e+17, 1.291629523605078e+17, 1.291629523637892e+17, 1.291629523669142e+17, 1.291629523701953e+17, 1.291629523733203e+17, 1.291629523766016e+17, 1.291629523798829e+17, 1.291629523830079e+17, 1.291629523862892e+17, 1.291629523894141e+17, 1.291629523926953e+17, 1.291629523959766e+17, 1.291629523991017e+17, 1.291629524023828e+17, 1.291629524056641e+17, 1.291629524087891e+17, 1.291629524120704e+17, 1.291629524151953e+17, 1.291629524184767e+17, 1.291629524216017e+17, 1.291629524248828e+17, 1.291629524281641e+17, 1.291629524312892e+17, 1.291629524345704e+17, 1.291629524376954e+17, 1.291629524409766e+17, 1.291629524442579e+17, 1.291629524473828e+17, 1.291629524506642e+17, 1.291629524539453e+17, 1.291629524570703e+17, 1.291629524603516e+17, 1.291629524634766e+17, 1.291629524667579e+17, 1.291629524698828e+17, 1.291629524731642e+17, 1.291629524764453e+17, 1.291629524795703e+17, 1.291629524828516e+17, 1.291629524859767e+17, 1.291629524892579e+17, 1.291629524925391e+17, 1.291629524956641e+17, 1.291629524989454e+17, 1.291629525020703e+17, 1.291629525053517e+17, 1.291629525086328e+17, 1.291629525117578e+17, 1.291629525150391e+17, 1.291629525181641e+17, 1.291629525214454e+17, 1.291629525247267e+17, 1.291629525278516e+17, 1.291629525311328e+17, 1.291629525342578e+17, 1.291629525375391e+17, 1.291629525408204e+17, 1.291629525439453e+17, 1.291629525472266e+17, 1.291629525503516e+17, 1.291629525536329e+17, 1.29162952556914e+17, 1.291629525600392e+17, 1.291629525633203e+17, 1.291629525666016e+17, 1.291629525697266e+17, 1.291629525730079e+17, 1.291629525761329e+17, 1.291629525794141e+17, 1.291629525826953e+17, 1.291629525858204e+17, 1.291629525891016e+17, 1.291629525922267e+17, 1.291629525955078e+17, 1.291629525987891e+17, 1.291629526019141e+17, 1.291629526051954e+17, 1.291629526083204e+17, 1.291629526116015e+17, 1.291629526148828e+17, 1.291629526181641e+17, 1.291629526212891e+17, 1.291629526245704e+17, 1.291629526276954e+17, 1.291629526309765e+17, 1.291629526341016e+17, 1.291629526373828e+17, 1.291629526406641e+17, 1.291629526437891e+17, 1.291629526470703e+17, 1.291629526501953e+17, 1.291629526534766e+17, 1.291629526567579e+17, 1.291629526598829e+17, 1.29162952663164e+17, 1.291629526662892e+17, 1.291629526695703e+17, 1.291629526728516e+17, 1.291629526759766e+17, 1.291629526792579e+17, 1.291629526823828e+17, 1.291629526856641e+17, 1.291629526889454e+17, 1.291629526920704e+17, 1.291629526953516e+17, 1.291629526984765e+17, 1.291629527017578e+17, 1.291629527050391e+17, 1.291629527081641e+17, 1.291629527114454e+17, 1.291629527145704e+17, 1.291629527178515e+17, 1.291629527211329e+17, 1.291629527242578e+17, 1.291629527275391e+17, 1.291629527306641e+17, 1.291629527339453e+17, 1.291629527372265e+17, 1.291629527403516e+17, 1.291629527436329e+17, 1.291629527467579e+17, 1.29162952750039e+17, 1.291629527533204e+17, 1.291629527564453e+17, 1.291629527597266e+17, 1.291629527630079e+17, 1.291629527661329e+17, 1.29162952769414e+17, 1.29162952772539e+17, 1.291629527758204e+17, 1.291629527791016e+17, 1.291629527822266e+17, 1.291629527855078e+17, 1.291629527886328e+17, 1.29162952791914e+17, 1.291629527951954e+17, 1.291629527983204e+17, 1.291629528016015e+17, 1.291629528047265e+17, 1.291629528080079e+17, 1.291629528112891e+17, 1.291629528144141e+17, 1.291629528176954e+17, 1.291629528208204e+17, 1.291629528241015e+17, 1.291629528273829e+17, 1.291629528305079e+17, 1.291629528337891e+17, 1.29162952836914e+17, 1.291629528401955e+17, 1.291629528434766e+17, 1.291629528466016e+17, 1.291629528498829e+17, 1.291629528530079e+17, 1.29162952856289e+17, 1.29162952859414e+17, 1.291629528626954e+17, 1.291629528659766e+17, 1.291629528691016e+17, 1.291629528723828e+17, 1.291629528756641e+17, 1.29162952878789e+17, 1.291629528820704e+17, 1.291629528851954e+17, 1.291629528884765e+17, 1.291629528917578e+17, 1.291629528948829e+17, 1.291629528981641e+17, 1.291629529012891e+17, 1.291629529045704e+17, 1.291629529076954e+17, 1.291629529109765e+17, 1.291629529142579e+17, 1.291629529173829e+17, 1.291629529206641e+17, 1.291629529237891e+17, 1.291629529270703e+17, 1.291629529303516e+17, 1.291629529334766e+17, 1.291629529367579e+17, 1.291629529398829e+17, 1.29162952943164e+17, 1.291629529464454e+17, 1.291629529495704e+17, 1.291629529528516e+17, 1.291629529559766e+17, 1.291629529592579e+17, 1.291629529625391e+17, 1.29162952965664e+17, 1.291629529689454e+17, 1.291629529720704e+17, 1.291629529753516e+17, 1.291629529786328e+17, 1.29162952981758e+17, 1.291629529850391e+17, 1.291629529881641e+17, 1.291629529914454e+17, 1.291629529947267e+17, 1.291629529978515e+17, 1.291629530011329e+17, 1.291629530044141e+17, 1.291629530075391e+17, 1.291629530108204e+17, 1.291629530139453e+17, 1.291629530172266e+17, 1.291629530205079e+17, 1.291629530236329e+17, 1.29162953026914e+17, 1.29162953030039e+17, 1.291629530333203e+17, 1.291629530366016e+17, 1.291629530397266e+17, 1.291629530430079e+17, 1.291629530461329e+17, 1.291629530494141e+17, 1.291629530526954e+17, 1.291629530558204e+17, 1.291629530591016e+17, 1.291629530623828e+17, 1.291629530655078e+17, 1.291629530687891e+17, 1.291629530719141e+17, 1.291629530751954e+17, 1.291629530784765e+17, 1.291629530816015e+17, 1.291629530848828e+17, 1.291629530880079e+17, 1.291629530912891e+17, 1.291629530945704e+17, 1.291629530976954e+17, 1.291629531009766e+17, 1.291629531041016e+17, 1.291629531073829e+17, 1.291629531106641e+17, 1.291629531137891e+17, 1.291629531170703e+17, 1.291629531201953e+17, 1.291629531234766e+17, 1.291629531267579e+17, 1.291629531298829e+17, 1.29162953133164e+17, 1.291629531362892e+17, 1.291629531395704e+17, 1.291629531428516e+17, 1.291629531459766e+17, 1.291629531492579e+17, 1.291629531523828e+17, 1.291629531556641e+17, 1.291629531589453e+17, 1.291629531620704e+17, 1.291629531653516e+17, 1.291629531684765e+17, 1.291629531717578e+17, 1.291629531750391e+17, 1.291629531781641e+17, 1.291629531814454e+17, 1.291629531847267e+17, 1.291629531878515e+17, 1.291629531911328e+17, 1.291629531942579e+17, 1.291629531975391e+17, 1.291629532006641e+17, 1.291629532039453e+17, 1.291629532072266e+17, 1.291629532103516e+17, 1.291629532136329e+17, 1.291629532167579e+17, 1.29162953220039e+17, 1.291629532233203e+17, 1.291629532264454e+17, 1.291629532297266e+17, 1.291629532328516e+17, 1.291629532361329e+17, 1.291629532394141e+17, 1.291629532425391e+17, 1.291629532458203e+17, 1.291629532491017e+17, 1.291629532522266e+17, 1.291629532555078e+17, 1.291629532586328e+17, 1.291629532619141e+17, 1.291629532651953e+17, 1.291629532683204e+17, 1.291629532716017e+17, 1.291629532747265e+17, 1.291629532780078e+17, 1.291629532812891e+17, 1.291629532844141e+17, 1.291629532876954e+17, 1.291629532908204e+17, 1.291629532941016e+17, 1.291629532973828e+17, 1.291629533005078e+17, 1.291629533037892e+17, 1.29162953306914e+17, 1.291629533101953e+17, 1.291629533134766e+17, 1.291629533166016e+17, 1.291629533198828e+17, 1.291629533230079e+17, 1.291629533262892e+17, 1.29162953329414e+17, 1.291629533326953e+17, 1.291629533359766e+17, 1.291629533391016e+17, 1.291629533423828e+17, 1.291629533456641e+17, 1.291629533487891e+17, 1.291629533520703e+17, 1.291629533551954e+17, 1.291629533584767e+17, 1.291629533617578e+17, 1.291629533648828e+17, 1.291629533681641e+17, 1.291629533712891e+17, 1.291629533745702e+17, 1.291629533778516e+17, 1.291629533809766e+17, 1.291629533842578e+17, 1.291629533873828e+17, 1.291629533906642e+17, 1.291629533939453e+17, 1.291629533970703e+17, 1.291629534003516e+17, 1.291629534036329e+17, 1.291629534067578e+17, 1.291629534100392e+17, 1.291629534131642e+17, 1.291629534164453e+17, 1.291629534197266e+17, 1.291629534228516e+17, 1.291629534261329e+17, 1.291629534292579e+17, 1.291629534325391e+17, 1.291629534358203e+17, 1.291629534389453e+17, 1.291629534422266e+17, 1.291629534453517e+17, 1.291629534486328e+17, 1.291629534519141e+17, 1.291629534550391e+17, 1.291629534583204e+17, 1.291629534614452e+17, 1.291629534647267e+17, 1.291629534680078e+17, 1.291629534711328e+17, 1.291629534744141e+17, 1.291629534776954e+17, 1.291629534808204e+17, 1.291629534841016e+17, 1.291629534872266e+17, 1.291629534905078e+17, 1.291629534937892e+17, 1.291629534969142e+17, 1.291629535001953e+17, 1.291629535033203e+17, 1.291629535066016e+17, 1.291629535098829e+17, 1.291629535130079e+17, 1.291629535162892e+17, 1.291629535194141e+17, 1.291629535226953e+17, 1.291629535259767e+17, 1.291629535291016e+17, 1.291629535323828e+17, 1.291629535355078e+17, 1.291629535387891e+17, 1.291629535420703e+17, 1.291629535451954e+17, 1.291629535484767e+17, 1.291629535516017e+17, 1.291629535548828e+17, 1.291629535581641e+17, 1.291629535612891e+17, 1.291629535645704e+17, 1.291629535676954e+17, 1.291629535709766e+17, 1.291629535742578e+17, 1.291629535773828e+17, 1.291629535806642e+17, 1.291629535837891e+17, 1.291629535870703e+17, 1.291629535903516e+17, 1.291629535934766e+17, 1.291629535967578e+17, 1.291629535998829e+17, 1.291629536031642e+17, 1.291629536064453e+17, 1.291629536095703e+17, 1.291629536128517e+17, 1.291629536159766e+17, 1.291629536192579e+17, 1.291629536223828e+17, 1.291629536256641e+17, 1.291629536289453e+17, 1.291629536322266e+17, 1.291629536353517e+17, 1.291629536386328e+17, 1.291629536417578e+17, 1.291629536450391e+17, 1.291629536483204e+17, 1.291629536514454e+17, 1.291629536547267e+17, 1.291629536580079e+17, 1.291629536611328e+17, 1.291629536644141e+17, 1.291629536675392e+17, 1.291629536708204e+17, 1.291629536739453e+17, 1.291629536772266e+17, 1.291629536805079e+17, 1.291629536836328e+17, 1.291629536869142e+17, 1.291629536901953e+17, 1.291629536933203e+17, 1.291629536966016e+17, 1.291629536997267e+17, 1.291629537030079e+17, 1.29162953706289e+17, 1.291629537094141e+17, 1.291629537126954e+17, 1.291629537158203e+17, 1.291629537191016e+17, 1.291629537223828e+17, 1.291629537255078e+17, 1.291629537287891e+17, 1.291629537319141e+17, 1.291629537351954e+17, 1.291629537384765e+17, 1.291629537416017e+17, 1.291629537448828e+17, 1.291629537480078e+17, 1.291629537512891e+17, 1.291629537545704e+17, 1.291629537576954e+17, 1.291629537609765e+17, 1.291629537641016e+17, 1.291629537673829e+17, 1.291629537706641e+17, 1.291629537737891e+17, 1.291629537770703e+17, 1.291629537801953e+17, 1.291629537834766e+17, 1.291629537867579e+17, 1.291629537898829e+17, 1.29162953793164e+17, 1.291629537962892e+17, 1.291629537995704e+17, 1.291629538028516e+17, 1.291629538059766e+17, 1.291629538092579e+17, 1.291629538123828e+17, 1.291629538156641e+17, 1.291629538189454e+17, 1.291629538220704e+17, 1.291629538253516e+17, 1.291629538284767e+17, 1.291629538317578e+17, 1.291629538348828e+17, 1.291629538381641e+17, 1.291629538414454e+17, 1.291629538445704e+17, 1.291629538478515e+17, 1.291629538511328e+17, 1.291629538542579e+17, 1.291629538575391e+17, 1.291629538606641e+17, 1.291629538639453e+17, 1.291629538672266e+17, 1.291629538703516e+17, 1.291629538736329e+17, 1.291629538767579e+17, 1.29162953880039e+17, 1.291629538831642e+17, 1.291629538864453e+17, 1.291629538897266e+17, 1.291629538928516e+17, 1.291629538961329e+17, 1.291629538992579e+17, 1.291629539025391e+17, 1.291629539058204e+17, 1.291629539089454e+17, 1.291629539122266e+17, 1.291629539153517e+17, 1.291629539186328e+17, 1.291629539219141e+17, 1.291629539250391e+17, 1.291629539283204e+17, 1.291629539316015e+17, 1.291629539347265e+17, 1.291629539380078e+17, 1.291629539411329e+17, 1.291629539444141e+17, 1.291629539476954e+17, 1.291629539508204e+17, 1.291629539541016e+17, 1.291629539572266e+17, 1.291629539605079e+17, 1.291629539637891e+17, 1.29162953966914e+17, 1.291629539701953e+17, 1.291629539734766e+17, 1.291629539766016e+17, 1.291629539798829e+17, 1.29162953983164e+17, 1.29162953986289e+17, 1.291629539895704e+17, 1.291629539926953e+17, 1.291629539959766e+17, 1.291629539992579e+17, 1.291629540023828e+17, 1.29162954005664e+17, 1.291629540087891e+17, 1.291629540120704e+17, 1.291629540151954e+17, 1.291629540184765e+17, 1.29162954021758e+17, 1.291629540248828e+17, 1.291629540281641e+17, 1.291629540314454e+17, 1.291629540345704e+17, 1.291629540378515e+17, 1.291629540409765e+17, 1.291629540442579e+17, 1.291629540475391e+17, 1.291629540506641e+17, 1.291629540539453e+17, 1.291629540570703e+17, 1.291629540603516e+17, 1.291629540636329e+17, 1.291629540667579e+17, 1.29162954070039e+17, 1.29162954073164e+17, 1.291629540764454e+17, 1.291629540797266e+17, 1.291629540828516e+17, 1.291629540861329e+17, 1.291629540892579e+17, 1.29162954092539e+17, 1.291629540958204e+17, 1.291629540989454e+17, 1.291629541022266e+17, 1.291629541053516e+17, 1.29162954108633e+17, 1.291629541119141e+17, 1.291629541150391e+17, 1.291629541183204e+17, 1.291629541214454e+17, 1.291629541247265e+17, 1.291629541280079e+17, 1.291629541311329e+17, 1.291629541344141e+17, 1.291629541375391e+17, 1.291629541408204e+17, 1.291629541441016e+17, 1.291629541472265e+17, 1.291629541505079e+17, 1.291629541536329e+17, 1.29162954156914e+17, 1.291629541601953e+17, 1.291629541633204e+17, 1.291629541666016e+17, 1.291629541697266e+17, 1.291629541730079e+17, 1.291629541762892e+17, 1.29162954179414e+17, 1.291629541826954e+17, 1.291629541858204e+17, 1.291629541891016e+17, 1.291629541923828e+17, 1.291629541955078e+17, 1.291629541987891e+17, 1.291629542019141e+17, 1.291629542051954e+17, 1.291629542084767e+17, 1.291629542116015e+17, 1.291629542148829e+17, 1.291629542180079e+17, 1.291629542212891e+17, 1.291629542244141e+17, 1.291629542276954e+17, 1.291629542309766e+17, 1.291629542341015e+17, 1.291629542373829e+17, 1.291629542405079e+17, 1.291629542437891e+17, 1.291629542470703e+17, 1.291629542501955e+17, 1.291629542534766e+17, 1.291629542566016e+17, 1.291629542598829e+17, 1.291629542631642e+17, 1.29162954266289e+17, 1.291629542695704e+17, 1.291629542728516e+17, 1.291629542759766e+17, 1.291629542792579e+17, 1.291629542823828e+17, 1.291629542856641e+17, 1.291629542889454e+17, 1.291629542920704e+17, 1.291629542953516e+17, 1.291629542984765e+17, 1.291629543017578e+17, 1.291629543048829e+17, 1.291629543081641e+17, 1.291629543114454e+17, 1.291629543147265e+17, 1.291629543178516e+17, 1.291629543211328e+17, 1.291629543242579e+17, 1.291629543275391e+17, 1.291629543308204e+17, 1.291629543339453e+17, 1.291629543372266e+17, 1.291629543405078e+17, 1.291629543436329e+17, 1.29162954346914e+17, 1.291629543500392e+17, 1.291629543533203e+17, 1.291629543564454e+17, 1.291629543597266e+17, 1.291629543630079e+17, 1.291629543661329e+17, 1.291629543694141e+17, 1.291629543726953e+17, 1.291629543758204e+17, 1.291629543791016e+17, 1.291629543822266e+17, 1.291629543855078e+17, 1.291629543886328e+17, 1.291629543919141e+17, 1.291629543951953e+17, 1.291629543983204e+17, 1.291629544016015e+17, 1.291629544048828e+17, 1.291629544080078e+17, 1.291629544112891e+17, 1.291629544144141e+17, 1.291629544176954e+17, 1.291629544209766e+17, 1.291629544241016e+17, 1.291629544273828e+17, 1.291629544305079e+17, 1.291629544337891e+17, 1.291629544370703e+17, 1.291629544401953e+17, 1.291629544434766e+17, 1.291629544466016e+17, 1.291629544498829e+17, 1.291629544531642e+17, 1.29162954456289e+17, 1.291629544595703e+17, 1.291629544626954e+17, 1.291629544659766e+17, 1.291629544692579e+17, 1.291629544723828e+17, 1.291629544756641e+17, 1.291629544787891e+17, 1.291629544820703e+17, 1.291629544853517e+17, 1.291629544884765e+17, 1.291629544917578e+17, 1.291629544948828e+17, 1.291629544981641e+17, 1.291629545014452e+17, 1.291629545045704e+17, 1.291629545078516e+17, 1.291629545109766e+17, 1.291629545142578e+17, 1.291629545175392e+17, 1.291629545206641e+17, 1.291629545239453e+17, 1.291629545270703e+17, 1.291629545303516e+17, 1.291629545336328e+17, 1.291629545367578e+17, 1.291629545400392e+17, 1.29162954543164e+17, 1.291629545464453e+17, 1.291629545497266e+17, 1.291629545528516e+17, 1.291629545561327e+17, 1.291629545592579e+17, 1.291629545625391e+17, 1.291629545658203e+17, 1.291629545689453e+17, 1.291629545722267e+17, 1.291629545753516e+17, 1.291629545786328e+17, 1.291629545819141e+17, 1.291629545850391e+17, 1.291629545883203e+17, 1.291629545914454e+17, 1.291629545947267e+17, 1.291629545980078e+17, 1.291629546011328e+17, 1.291629546044141e+17, 1.291629546075391e+17, 1.291629546108204e+17, 1.291629546141016e+17, 1.291629546172266e+17, 1.291629546205078e+17, 1.291629546236328e+17, 1.291629546269142e+17, 1.291629546301953e+17, 1.291629546333203e+17, 1.291629546366016e+17, 1.291629546398829e+17, 1.291629546430077e+17, 1.291629546462892e+17, 1.291629546494141e+17, 1.291629546526953e+17, 1.291629546559766e+17, 1.291629546591017e+17, 1.291629546623828e+17, 1.291629546655078e+17, 1.291629546687891e+17, 1.291629546720704e+17, 1.291629546751953e+17, 1.291629546784767e+17, 1.291629546816017e+17, 1.291629546848828e+17, 1.291629546881641e+17, 1.291629546912891e+17, 1.291629546945704e+17, 1.291629546976952e+17, 1.291629547009766e+17, 1.291629547042578e+17, 1.291629547073828e+17, 1.291629547106641e+17, 1.291629547137892e+17, 1.291629547170703e+17, 1.291629547203516e+17, 1.291629547234766e+17, 1.291629547267579e+17, 1.291629547298828e+17, 1.291629547331642e+17, 1.291629547364453e+17, 1.291629547395703e+17, 1.291629547428516e+17, 1.291629547459766e+17, 1.291629547492579e+17, 1.291629547525391e+17, 1.291629547556641e+17, 1.291629547589454e+17, 1.291629547620703e+17, 1.291629547653517e+17, 1.291629547686328e+17, 1.291629547717578e+17, 1.291629547750391e+17, 1.291629547781641e+17, 1.291629547814454e+17, 1.291629547847267e+17, 1.291629547878516e+17, 1.291629547911328e+17, 1.291629547942578e+17, 1.291629547975391e+17, 1.291629548008204e+17, 1.291629548039453e+17, 1.291629548072266e+17, 1.291629548103516e+17, 1.291629548136329e+17, 1.291629548169142e+17, 1.291629548200392e+17, 1.291629548233203e+17, 1.291629548264453e+17, 1.291629548297266e+17, 1.291629548330079e+17, 1.291629548361329e+17, 1.291629548394141e+17, 1.291629548425391e+17, 1.291629548458203e+17, 1.291629548491017e+17, 1.291629548522266e+17, 1.291629548555078e+17, 1.291629548586328e+17, 1.291629548619141e+17, 1.291629548651953e+17, 1.291629548683204e+17, 1.291629548716017e+17, 1.291629548747267e+17, 1.291629548780078e+17, 1.291629548812891e+17, 1.291629548844141e+17, 1.291629548876954e+17, 1.291629548908204e+17, 1.291629548941016e+17, 1.291629548973828e+17, 1.291629549005079e+17, 1.291629549037892e+17, 1.291629549069142e+17, 1.291629549101953e+17, 1.291629549134766e+17, 1.291629549166016e+17, 1.291629549198829e+17, 1.29162954923164e+17, 1.291629549262892e+17, 1.291629549295703e+17, 1.291629549326953e+17, 1.291629549359766e+17, 1.291629549392579e+17, 1.291629549423828e+17, 1.291629549456641e+17, 1.291629549487891e+17, 1.291629549520703e+17, 1.291629549553516e+17, 1.291629549584767e+17, 1.291629549617578e+17, 1.291629549648828e+17, 1.291629549681641e+17, 1.291629549714454e+17, 1.291629549745704e+17, 1.291629549778516e+17, 1.291629549809766e+17, 1.291629549842578e+17, 1.291629549873828e+17, 1.291629549906642e+17, 1.291629549939453e+17, 1.291629549970703e+17, 1.291629550003516e+17, 1.291629550036329e+17, 1.291629550067578e+17, 1.29162955010039e+17, 1.291629550133203e+17, 1.291629550164453e+17, 1.291629550197266e+17, 1.291629550228516e+17, 1.291629550261329e+17, 1.29162955029414e+17, 1.291629550325391e+17, 1.291629550358204e+17, 1.291629550389453e+17, 1.291629550422266e+17, 1.291629550455078e+17, 1.291629550486328e+17, 1.291629550519141e+17, 1.291629550550391e+17, 1.291629550583204e+17, 1.291629550616015e+17, 1.291629550647267e+17, 1.291629550680079e+17, 1.291629550711328e+17, 1.291629550744141e+17, 1.291629550776954e+17, 1.291629550808204e+17, 1.291629550841015e+17, 1.291629550872266e+17, 1.291629550905079e+17, 1.291629550937891e+17, 1.29162955096914e+17, 1.291629551001953e+17, 1.291629551033203e+17, 1.291629551066016e+17, 1.291629551098829e+17, 1.291629551130079e+17, 1.29162955116289e+17, 1.291629551194141e+17, 1.291629551226954e+17, 1.291629551259766e+17, 1.291629551291016e+17, 1.291629551323828e+17, 1.291629551355078e+17, 1.291629551387891e+17, 1.291629551420704e+17, 1.291629551451954e+17, 1.291629551484765e+17, 1.291629551516017e+17, 1.291629551548828e+17, 1.291629551581641e+17, 1.291629551612891e+17, 1.291629551645704e+17, 1.291629551676954e+17, 1.291629551709765e+17, 1.291629551742579e+17, 1.291629551773829e+17, 1.291629551806641e+17, 1.291629551839453e+17, 1.291629551870703e+17, 1.291629551903516e+17, 1.291629551934766e+17, 1.291629551967579e+17, 1.291629551998829e+17, 1.29162955203164e+17, 1.291629552064453e+17, 1.291629552095704e+17, 1.291629552128516e+17, 1.291629552161329e+17, 1.291629552192579e+17, 1.291629552225391e+17, 1.291629552256641e+17, 1.291629552289454e+17, 1.291629552320704e+17, 1.291629552353516e+17, 1.291629552386328e+17, 1.291629552417578e+17, 1.291629552450391e+17, 1.291629552481641e+17, 1.291629552514454e+17, 1.291629552547265e+17, 1.291629552578515e+17, 1.291629552611328e+17, 1.291629552642579e+17, 1.291629552675391e+17, 1.291629552708204e+17, 1.291629552739453e+17, 1.291629552772266e+17, 1.291629552805079e+17, 1.291629552836329e+17, 1.29162955286914e+17, 1.29162955290039e+17, 1.291629552933203e+17, 1.291629552964453e+17, 1.291629552997266e+17, 1.291629553030079e+17, 1.291629553061329e+17, 1.291629553094141e+17, 1.291629553126954e+17, 1.291629553158204e+17, 1.291629553191016e+17, 1.291629553222266e+17, 1.291629553255078e+17, 1.291629553286328e+17, 1.291629553319141e+17, 1.291629553351954e+17, 1.291629553383204e+17, 1.291629553416015e+17, 1.291629553448829e+17, 1.291629553480078e+17, 1.291629553512891e+17, 1.291629553545704e+17, 1.291629553576954e+17, 1.291629553609765e+17, 1.291629553641016e+17, 1.291629553673829e+17, 1.291629553706641e+17, 1.291629553737891e+17, 1.291629553770705e+17, 1.291629553801953e+17, 1.291629553834766e+17, 1.291629553867579e+17, 1.291629553898829e+17, 1.29162955393164e+17, 1.29162955396289e+17, 1.291629553995704e+17, 1.291629554028516e+17, 1.291629554059766e+17, 1.291629554092579e+17, 1.291629554123828e+17, 1.29162955415664e+17, 1.291629554189454e+17, 1.291629554220704e+17, 1.291629554253516e+17, 1.291629554284765e+17, 1.29162955431758e+17, 1.291629554350391e+17, 1.291629554381641e+17, 1.291629554414454e+17, 1.291629554445704e+17, 1.291629554478515e+17, 1.291629554511329e+17, 1.291629554542579e+17, 1.291629554575391e+17, 1.291629554606641e+17, 1.291629554639455e+17, 1.291629554672266e+17, 1.291629554703516e+17, 1.291629554736329e+17, 1.291629554767579e+17, 1.29162955480039e+17, 1.291629554833203e+17, 1.291629554864454e+17, 1.291629554897266e+17, 1.291629554928516e+17, 1.291629554961329e+17, 1.291629554994141e+17, 1.29162955502539e+17, 1.291629555058204e+17, 1.291629555089454e+17, 1.291629555122266e+17, 1.291629555155078e+17, 1.29162955518633e+17, 1.291629555219141e+17, 1.291629555250391e+17, 1.291629555283204e+17, 1.291629555316017e+17, 1.291629555347265e+17, 1.291629555380079e+17, 1.291629555411329e+17, 1.291629555444141e+17, 1.291629555476954e+17, 1.291629555508204e+17, 1.291629555541016e+17, 1.291629555573828e+17, 1.291629555605079e+17, 1.291629555637891e+17, 1.29162955566914e+17, 1.291629555701953e+17, 1.291629555733204e+17, 1.291629555766016e+17, 1.291629555798829e+17, 1.291629555830079e+17, 1.291629555862892e+17, 1.29162955589414e+17, 1.291629555926954e+17, 1.291629555959766e+17, 1.291629555991016e+17, 1.291629556023828e+17},
			             {1.291629441639453e+17, 1.291629441672266e+17, 1.291629441703516e+17, 1.291629441736329e+17, 1.29162944176914e+17, 1.291629441800392e+17, 1.291629441833203e+17, 1.291629441864453e+17, 1.291629441897266e+17, 1.291629441928516e+17, 1.291629441961329e+17, 1.29162944199414e+17, 1.291629442025391e+17, 1.291629442058204e+17, 1.291629442089453e+17, 1.291629442122266e+17, 1.291629442155078e+17, 1.291629442186328e+17, 1.291629442219141e+17, 1.291629442250391e+17, 1.291629442283204e+17, 1.291629442316015e+17, 1.291629442347267e+17, 1.291629442380079e+17, 1.291629442411328e+17, 1.291629442444141e+17, 1.291629442476954e+17, 1.291629442508204e+17, 1.291629442541015e+17, 1.291629442572266e+17, 1.291629442605079e+17, 1.291629442636328e+17, 1.29162944266914e+17, 1.291629442701953e+17, 1.291629442733203e+17, 1.291629442766016e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
