netcdf mask {
	:date_created = "20200811T114915";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200811T114915";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 28;
			channels = 6;
			categories = 168;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  77.9, 79.2, 64.6, 79.0, 73.3, 80.1, 81.1, 46.5, 76.3, 74.8, 73.5, 79.0, 78.8, 79.0, 80.4, 76.5, 74.5, 79.6, 80.0, 79.7, 78.0, 79.9, 80.4, 72.4, 73.9, 78.7, 79.0, 79.5;
			max_depth =  80.5, 80.9, 78.7, 81.4, 82.0, 81.5, 82.7, 53.7, 83.1, 77.7, 75.3, 81.1, 81.2, 80.7, 81.5, 78.2, 76.2, 81.0, 81.1, 81.1, 79.5, 81.1, 80.9, 73.6, 76.3, 80.0, 80.9, 80.8;
			start_time = 130432232097982080, 130432232251888256, 130432233157357056, 130432233727513216, 130432234533607040, 130432233935638272, 130432235800481920, 130432254258919424, 130432256195481984, 130432268758294528, 130432270831263232, 130432268648919424, 130432268890950784, 130432237320794496, 130432261229232000, 130432261568919552, 130432261938606976, 130432263681575808, 130432264761107072, 130432264938606976, 130432264945794432, 130432265286107008, 130432263955950720, 130432267766575744, 130432267855481984, 130432270270482048, 130432275282356992, 130432275845638272;
			end_time = 130432232143294464, 130432232342513152, 130432233220482048, 130432233772825728, 130432234597044480, 130432233971888256, 130432235827669504, 130432254421731968, 130432256313138304, 130432268913450752, 130432270941575680, 130432268802513152, 130432269031263360, 130432237347825792, 130432261258919552, 130432261605950720, 130432262012513152, 130432263822669568, 130432264909075712, 130432265042044416, 130432265034388352, 130432265367200768, 130432264029388160, 130432267907044480, 130432267959075712, 130432270345325824, 130432275380169472, 130432275913607040;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21","Layer22","Layer23","Layer24","Layer25","Layer26","Layer27","Layer28";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "6007", "6007", "6007", "6007", "6007", "6007", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "6007", "6007", "6007", "6007", "6007", "6007", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "6007", "6007", "6007", "6007", "6007", "6007", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63;
			mask_times = {1.304322320979821e+17, 1.304322321070445e+17, 1.30432232116107e+17, 1.304322321251695e+17, 1.304322321432945e+17},
			             {1.304322322518883e+17, 1.304322322609508e+17, 1.304322322700133e+17, 1.304322322790757e+17, 1.304322322881382e+17, 1.304322322972008e+17, 1.304322323062633e+17, 1.30432232315482e+17, 1.304322323243882e+17, 1.304322323334508e+17, 1.304322323425132e+17},
			             {1.304322331573571e+17, 1.304322331664196e+17, 1.304322331753257e+17, 1.30432233220482e+17},
			             {1.304322337275132e+17, 1.304322337365757e+17, 1.304322337454821e+17, 1.304322337545445e+17, 1.304322337637632e+17, 1.304322337728257e+17},
			             {1.30432234533607e+17, 1.304322345426694e+17, 1.304322345518883e+17, 1.304322345607945e+17, 1.304322345879821e+17, 1.304322345970445e+17},
			             {1.304322339356383e+17, 1.304322339718883e+17},
			             {1.304322358004819e+17, 1.304322358095444e+17, 1.304322358276695e+17},
			             {1.304322542589194e+17, 1.30432254421732e+17},
			             {1.30432256195482e+17, 1.304322562045445e+17, 1.304322562317321e+17, 1.304322562407945e+17, 1.30432256249857e+17, 1.304322562589196e+17, 1.30432256267982e+17, 1.304322562770445e+17, 1.30432256286107e+17, 1.304322563040758e+17, 1.304322563131383e+17},
			             {1.304322687582945e+17, 1.304322687659507e+17, 1.30432268772982e+17, 1.304322687803258e+17, 1.304322688097007e+17, 1.304322688170445e+17, 1.304322688318883e+17, 1.30432268839232e+17, 1.304322688465757e+17, 1.304322688540758e+17, 1.304322688837632e+17, 1.304322688909508e+17, 1.304322688987633e+17, 1.30432268906107e+17, 1.304322689134508e+17},
			             {1.304322708312632e+17, 1.304322708678258e+17, 1.304322708751695e+17, 1.304322708825133e+17, 1.304322709048571e+17, 1.304322709120445e+17, 1.304322709193883e+17, 1.304322709415757e+17},
			             {1.304322686489194e+17, 1.304322686562633e+17, 1.30432268663607e+17, 1.304322686709508e+17, 1.304322686781382e+17, 1.30432268685482e+17, 1.304322686928257e+17, 1.304322687000133e+17, 1.304322687073571e+17, 1.304322687147008e+17, 1.304322687220445e+17, 1.30432268772982e+17, 1.304322687803258e+17, 1.304322687875132e+17, 1.304322687951695e+17, 1.304322688025132e+17},
			             {1.304322688909508e+17, 1.304322688987633e+17, 1.30432268906107e+17, 1.304322689134508e+17, 1.304322689207945e+17, 1.304322689281382e+17, 1.304322689353258e+17, 1.304322689428257e+17, 1.304322689501695e+17, 1.304322689576695e+17, 1.304322690020445e+17, 1.30432269009232e+17, 1.304322690165757e+17, 1.304322690239196e+17, 1.304322690312634e+17},
			             {1.304322373207945e+17, 1.304322373478258e+17},
			             {1.30432261229232e+17, 1.304322612589196e+17},
			             {1.304322615689196e+17, 1.304322616059507e+17},
			             {1.30432261938607e+17, 1.304322620125132e+17},
			             {1.304322636815758e+17, 1.304322636890757e+17, 1.304322637111069e+17, 1.30432263718607e+17, 1.30432263741732e+17, 1.304322637490757e+17, 1.304322637564195e+17, 1.304322637637632e+17, 1.304322637712632e+17, 1.304322637931382e+17, 1.30432263800482e+17, 1.304322638079821e+17, 1.304322638153257e+17, 1.304322638226696e+17},
			             {1.304322647611071e+17, 1.304322649090757e+17},
			             {1.30432264938607e+17, 1.304322650420444e+17},
			             {1.304322649457944e+17, 1.304322650343884e+17},
			             {1.30432265286107e+17, 1.304322653598569e+17, 1.304322653672008e+17},
			             {1.304322639559507e+17, 1.304322640293882e+17},
			             {1.304322677665757e+17, 1.304322679070445e+17},
			             {1.30432267855482e+17, 1.304322679590757e+17},
			             {1.30432270270482e+17, 1.304322703228257e+17, 1.304322703301696e+17, 1.304322703376695e+17, 1.304322703453258e+17},
			             {1.30432275282357e+17, 1.304322753131383e+17, 1.304322753211069e+17, 1.304322753801695e+17},
			             {1.304322758456383e+17, 1.304322758531382e+17, 1.304322758603258e+17, 1.304322758681382e+17, 1.304322758753258e+17, 1.304322758826696e+17, 1.304322758900133e+17, 1.30432275898607e+17, 1.30432275913607e+17};
			mask_depths = {{77.9, 80.4}, {77.9, 80.4}, {78.0, 80.5}, {77.9, 80.4}, {77.9, 80.4}}, {{79.2, 80.9}, {79.3}, {79.2}, {80.9}, {79.2, 80.8}, {79.3, 80.7, 80.9}, {79.2}, {80.5}, {79.2}, {79.3, 80.5}, {79.2, 80.4}}, {{64.6, 72.5}, {72.6, 72.7}, {72.8, 78.7}, {64.6, 78.7}}, {{79.0, 80.8}, {79.1, 80.8}, {79.0, 80.7}, {79.1, 80.8, 81.0}, {79.0, 81.1, 81.2}, {79.1, 81.3, 81.4}}, {{73.3, 81.9}, {81.8}, {81.8}, {81.9}, {73.3, 81.9}, {73.4, 82.0}}, {{80.1, 81.5}, {80.1, 81.5}}, {{81.1, 82.7}, {82.6}, {81.1, 82.6}}, {{46.5, 53.7}, {46.5, 53.7}}, {{76.4, 82.8}, {76.3, 82.9}, {76.3, 82.9}, {76.4}, {83.1}, {83.1}, {76.4, 83.0}, {76.5, 83.1}, {76.4, 83.1}, {82.9}, {76.4, 82.9}}, {{75.3, 77.7}, {75.3, 77.7}, {75.2, 77.6}, {75.3, 77.7}, {75.3, 77.7}, {75.2, 77.6}, {75.2, 77.6}, {75.3, 77.7}, {75.3, 77.7}, {75.2, 77.6}, {75.2, 77.6}, {75.3, 77.7}, {75.3, 77.3, 77.7}, {74.8, 75.1, 75.2, 77.2}, {75.2, 77.3, 77.6}}, {{73.5, 75.2}, {75.2}, {75.3}, {75.2}, {73.5, 75.2}, {73.6, 75.3}, {73.5, 75.2}, {73.5, 75.2}}, {{79.1, 80.3}, {79.1, 80.3}, {79.0, 80.2}, {80.3, 80.4}, {80.5, 80.7}, {79.0, 80.8}, {79.1}, {79.0}, {79.1}, {79.1, 80.8}, {79.0, 80.9}, {80.9}, {81.0}, {81.0}, {81.1}, {79.0, 81.1}}, {{79.3, 81.2}, {80.7, 81.1}, {78.8, 79.0, 79.1, 80.6}, {79.1, 80.7, 81.0}, {80.9}, {79.1}, {79.2, 80.9}, {79.2, 81.0}, {79.3, 81.0}, {79.2, 80.9}, {79.2}, {79.3}, {80.9}, {80.8}, {79.3, 80.8}}, {{79.0, 80.7}, {79.0, 80.7}}, {{80.4, 81.5}, {80.4, 81.5}}, {{76.5, 78.2}, {76.5, 78.2}}, {{74.5, 76.2}, {74.5, 76.2}}, {{79.6, 80.7}, {80.7}, {80.9, 81.0}, {80.8}, {80.8}, {80.9}, {80.8}, {80.8}, {80.9}, {80.9}, {81.0}, {80.9}, {80.9}, {79.6, 81.0}}, {{80.0, 81.1}, {80.0, 81.1}}, {{79.7, 81.1}, {79.7, 81.1}}, {{78.0, 79.5}, {78.0, 79.5}}, {{79.9, 81.0}, {81.0}, {79.9, 81.1}}, {{80.4, 80.9}, {80.4, 80.9}}, {{72.4, 73.6}, {72.4, 73.6}}, {{73.9, 76.3}, {73.9, 76.3}}, {{78.7, 79.9}, {79.9}, {80.0}, {79.9}, {78.7, 79.9}}, {{79.0, 80.8}, {80.8}, {80.9}, {79.0, 80.9}}, {{79.5, 80.7}, {80.7, 80.8}, {80.6}, {80.7}, {80.7}, {80.6}, {80.7}, {80.6}, {79.5, 80.6}};
		}
	}
}
