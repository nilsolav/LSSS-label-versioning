netcdf mask {
	:date_created = "20200810T140900";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200810T140900";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 28;
			channels = 6;
			categories = 168;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0, 15.0, 45.2, 32.9, 40.3, 49.1, 47.4, 49.1, 41.2, 51.7, 48.1, 49.2, 51.6, 45.7, 47.8, 49.9, 52.3, 46.4, 52.2, 55.9, 50.8, 49.7, 58.5, 55.5, 59.4, 53.6, 48.3, 51.9;
			max_depth =  61.7, 60.9, 50.0, 35.8, 44.2, 51.7, 52.1, 59.4, 48.3, 57.8, 55.2, 53.3, 54.6, 52.9, 50.7, 52.8, 56.0, 52.0, 55.9, 58.1, 55.7, 53.6, 60.3, 58.8, 61.4, 58.7, 58.3, 55.8;
			start_time = 131067417153558016, 131067433006526720, 131067418008401792, 131067417557308032, 131067418354339200, 131067418470745600, 131067430519964288, 131067430641526784, 131067427534495488, 131067427530276736, 131067427643714304, 131067427949182976, 131067422176683008, 131067423114339200, 131067419683870592, 131067424200901760, 131067425734964224, 131067426061839232, 131067431004495488, 131067431392464256, 131067431426683008, 131067431647620480, 131067431685745536, 131067424816214272, 131067432272464256, 131067432331995392, 131067432507776768, 131067432957151744;
			end_time = 131067433006526720, 131067439410276736, 131067418037620480, 131067417577464192, 131067418367620480, 131067418486995456, 131067430536214144, 131067430734339200, 131067427548089344, 131067427548089344, 131067427668558080, 131067427969964288, 131067422210120448, 131067423130901760, 131067419708401664, 131067424214026752, 131067425746995584, 131067426074339328, 131067431021995520, 131067431413245440, 131067431451526784, 131067431660120448, 131067431702464256, 131067424828401792, 131067432293870592, 131067432357151744, 131067432532151680, 131067432977933056;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28;
			region_name = "Layer1","Layer2","Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11","Layer12","Layer13","Layer14","Layer15","Layer16","Layer17","Layer18","Layer19","Layer20","Layer21","Layer22","Layer23","Layer24","Layer25","Layer26";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "27", "27", "27", "27", "27", "27", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010", "6010";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,   2,   3,   4,   5,   6,   7,   8,   9,  10,  11,  12,  13,  14,  15,  16,  17,  18,  19,  20,  21,  22,  23,  24,  25,  26,  27,  28,  29,  30,  31,  32,  33,  34,  35,  36,  37,  38,  39,  40,  41,  42,  43,  44,  45,  46,  47,  48,  49,  50,  51,  52,  53,  54,  55,  56,  57,  58,  59,  60,  61,  62,  63,  64,  65,  66,  67,  68,  69,  70,  71,  72,  73,  74,  75,  76,  77,  78,  79,  80,  81,  82,  83,  84,  85,  86,  87,  88,  89,  90,  91,  92,  93,  94,  95,  96,  97,  98,  99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63;
			mask_times = {1.31067417153558e+17, 1.310674171577768e+17, 1.310674171621518e+17, 1.31067417166058e+17, 1.310674171702767e+17, 1.310674171743393e+17, 1.310674171784017e+17, 1.310674171824643e+17, 1.310674171865268e+17, 1.310674171909018e+17, 1.310674171951205e+17, 1.310674171991831e+17, 1.31067417203558e+17, 1.310674172079331e+17, 1.31067417212308e+17, 1.310674172163706e+17, 1.31067417220433e+17, 1.310674172249642e+17, 1.310674172290268e+17, 1.31067417232933e+17, 1.310674172374643e+17, 1.310674172413705e+17, 1.310674172454331e+17, 1.310674172502769e+17, 1.310674172546518e+17, 1.310674172588705e+17, 1.31067417262933e+17, 1.310674172671517e+17, 1.310674172716831e+17, 1.310674172757455e+17, 1.31067417279808e+17, 1.31067417284183e+17, 1.310674172887142e+17, 1.310674172927768e+17, 1.31067417297308e+17, 1.310674173013705e+17, 1.31067417305433e+17, 1.310674173094956e+17, 1.310674173140269e+17, 1.310674173180892e+17, 1.31067417322308e+17, 1.310674173265267e+17, 1.310674173307455e+17, 1.310674173348081e+17, 1.31067417339183e+17, 1.310674173432456e+17, 1.31067417347308e+17, 1.310674173519955e+17, 1.31067417356058e+17, 1.310674173601206e+17, 1.310674173643392e+17, 1.310674173684017e+17, 1.31067417372933e+17, 1.31067417377308e+17, 1.310674173815268e+17, 1.310674173855892e+17, 1.310674173896517e+17, 1.310674173940268e+17, 1.310674173985581e+17, 1.310674174024643e+17, 1.310674174065268e+17, 1.310674174110579e+17, 1.310674174154331e+17, 1.310674174196517e+17, 1.310674174238705e+17, 1.310674174279331e+17, 1.310674174321517e+17, 1.310674174363704e+17, 1.310674174405892e+17, 1.310674174446518e+17, 1.310674174488705e+17, 1.31067417452933e+17, 1.310674174569955e+17, 1.310674174612143e+17, 1.310674174652768e+17, 1.310674174693393e+17, 1.310674174734017e+17, 1.310674174776205e+17, 1.310674174816831e+17, 1.310674174857454e+17, 1.31067417489808e+17, 1.310674174940268e+17, 1.310674174980893e+17, 1.310674175021517e+17, 1.310674175063704e+17, 1.310674175105892e+17, 1.310674175146518e+17, 1.310674175188705e+17, 1.310674175234017e+17, 1.310674175276205e+17, 1.310674175321518e+17, 1.310674175362143e+17, 1.310674175402767e+17, 1.310674175451205e+17, 1.310674175491831e+17, 1.310674175532454e+17, 1.31067417557308e+17, 1.310674175613705e+17, 1.310674175652767e+17, 1.310674175694956e+17, 1.310674175734019e+17, 1.310674175774642e+17, 1.310674175815268e+17, 1.310674175855892e+17, 1.31067417589808e+17, 1.310674175938705e+17, 1.310674175979331e+17, 1.310674176019955e+17, 1.310674176062143e+17, 1.310674176102767e+17, 1.31067417614183e+17, 1.310674176182455e+17, 1.310674176224643e+17, 1.310674176265267e+17, 1.310674176305893e+17, 1.310674176352767e+17, 1.310674176393393e+17, 1.310674176432456e+17, 1.310674176474643e+17, 1.310674176513705e+17, 1.310674176554331e+17, 1.310674176594954e+17, 1.31067417663558e+17, 1.310674176677768e+17, 1.310674176718392e+17, 1.31067417676058e+17, 1.310674176802767e+17, 1.310674176843392e+17, 1.310674176884018e+17, 1.310674176924643e+17, 1.310674176965267e+17, 1.310674177005892e+17, 1.310674177046518e+17, 1.310674177087142e+17, 1.310674177132456e+17, 1.31067417717308e+17, 1.310674177215267e+17, 1.310674177257455e+17, 1.31067417729808e+17, 1.31067417734183e+17, 1.310674177384017e+17, 1.310674177424643e+17, 1.31067417746683e+17, 1.310674177509018e+17, 1.310674177549642e+17, 1.310674177593393e+17, 1.31067417763558e+17, 1.310674177676205e+17, 1.310674177716829e+17, 1.310674177757455e+17, 1.310674177799643e+17, 1.310674177840268e+17, 1.310674177880892e+17, 1.31067417792308e+17, 1.310674177963706e+17, 1.310674178004329e+17, 1.310674178048081e+17, 1.310674178088704e+17, 1.31067417812933e+17, 1.31067417817308e+17, 1.310674178213705e+17, 1.310674178252767e+17, 1.310674178294956e+17, 1.31067417833558e+17, 1.310674178379331e+17, 1.310674178419955e+17, 1.310674178459017e+17, 1.310674178499643e+17, 1.310674178540268e+17, 1.310674178580892e+17, 1.310674178621518e+17, 1.310674178662143e+17, 1.310674178705893e+17, 1.310674178746518e+17, 1.310674178788705e+17, 1.310674178834017e+17, 1.310674178876205e+17, 1.310674178915268e+17, 1.310674178959017e+17, 1.310674178999643e+17, 1.310674179040268e+17, 1.310674179079329e+17, 1.310674179121517e+17, 1.310674179162143e+17, 1.310674179201204e+17, 1.31067417924183e+17, 1.310674179288705e+17, 1.31067417932933e+17, 1.310674179369955e+17, 1.31067417941058e+17, 1.310674179451205e+17, 1.31067417949183e+17, 1.310674179532456e+17, 1.310674179571517e+17, 1.310674179612142e+17, 1.310674179652768e+17, 1.310674179694956e+17, 1.310674179743393e+17, 1.310674179784017e+17, 1.310674179824643e+17, 1.31067417986683e+17, 1.310674179912142e+17, 1.310674179952768e+17, 1.310674179999643e+17, 1.310674180040268e+17, 1.310674180084018e+17, 1.310674180126205e+17, 1.31067418016683e+17, 1.310674180207455e+17, 1.310674180248081e+17, 1.310674180288704e+17, 1.31067418033558e+17, 1.310674180376205e+17, 1.310674180418392e+17, 1.310674180468393e+17, 1.310674180509018e+17, 1.310674180551205e+17, 1.310674180590268e+17, 1.310674180630893e+17, 1.310674180669955e+17, 1.310674180713705e+17, 1.31067418076058e+17, 1.310674180801204e+17, 1.310674180841829e+17, 1.310674180885581e+17, 1.310674180926204e+17, 1.310674180965267e+17, 1.310674181005892e+17, 1.310674181051205e+17, 1.31067418109183e+17, 1.310674181132454e+17, 1.31067418117308e+17, 1.310674181216831e+17, 1.310674181257455e+17, 1.31067418129808e+17, 1.310674181340268e+17, 1.310674181380892e+17, 1.310674181421517e+17, 1.310674181465267e+17, 1.310674181505893e+17, 1.310674181546516e+17, 1.310674181590268e+17, 1.31067418163558e+17, 1.310674181676205e+17, 1.310674181719955e+17, 1.31067418176058e+17, 1.310674181802767e+17, 1.310674181843392e+17, 1.310674181884017e+17, 1.310674181924643e+17, 1.310674181963704e+17, 1.310674182009018e+17, 1.310674182049642e+17, 1.310674182090268e+17, 1.310674182134017e+17, 1.310674182179331e+17, 1.310674182219955e+17, 1.310674182263704e+17, 1.31067418230433e+17, 1.310674182348079e+17, 1.310674182388705e+17, 1.310674182429331e+17, 1.310674182469955e+17, 1.310674182512142e+17, 1.310674182552768e+17, 1.310674182596517e+17, 1.310674182637143e+17, 1.310674182677768e+17, 1.310674182716831e+17, 1.310674182757455e+17, 1.31067418279808e+17, 1.310674182838705e+17, 1.310674182880892e+17, 1.31067418292308e+17, 1.310674182963706e+17, 1.310674183005893e+17, 1.310674183046516e+17, 1.310674183085581e+17, 1.310674183126204e+17, 1.31067418316683e+17, 1.310674183207456e+17, 1.310674183248079e+17, 1.310674183288704e+17, 1.310674183327768e+17, 1.310674183376205e+17, 1.310674183416829e+17, 1.310674183455894e+17, 1.310674183502767e+17, 1.310674183543392e+17, 1.310674183587142e+17, 1.310674183630893e+17, 1.310674183676205e+17, 1.310674183724643e+17, 1.310674183765268e+17, 1.310674183805892e+17, 1.310674183846518e+17, 1.310674183887142e+17, 1.310674183927767e+17, 1.31067418396683e+17, 1.310674184009018e+17, 1.310674184051205e+17, 1.31067418409183e+17, 1.310674184132456e+17, 1.31067418417308e+17, 1.310674184213705e+17, 1.310674184257455e+17, 1.31067418429808e+17, 1.310674184338705e+17, 1.310674184379331e+17, 1.310674184419955e+17, 1.310674184459018e+17, 1.310674184502767e+17, 1.310674184543393e+17, 1.310674184585581e+17, 1.310674184626204e+17, 1.31067418466683e+17, 1.310674184707456e+17, 1.310674184746518e+17, 1.310674184788704e+17, 1.31067418482933e+17, 1.310674184869955e+17, 1.310674184909018e+17, 1.310674184951205e+17, 1.310674184990267e+17, 1.310674185030893e+17, 1.310674185074642e+17, 1.310674185115268e+17, 1.310674185155892e+17, 1.310674185196517e+17, 1.310674185237143e+17, 1.310674185277768e+17, 1.310674185319955e+17, 1.310674185362143e+17, 1.310674185404329e+17, 1.310674185444955e+17, 1.310674185485581e+17, 1.310674185527768e+17, 1.310674185568392e+17, 1.310674185609018e+17, 1.310674185649644e+17, 1.310674185690267e+17, 1.310674185730893e+17, 1.31067418577308e+17, 1.310674185813705e+17, 1.31067418585433e+17, 1.310674185894954e+17, 1.31067418593558e+17, 1.310674185979329e+17, 1.310674186019955e+17, 1.310674186063704e+17, 1.31067418610433e+17, 1.310674186151205e+17, 1.310674186194956e+17, 1.310674186237143e+17, 1.310674186279329e+17, 1.310674186324643e+17, 1.310674186365268e+17, 1.310674186405892e+17, 1.310674186446518e+17, 1.310674186487142e+17, 1.310674186527767e+17, 1.310674186568393e+17, 1.310674186607455e+17, 1.310674186648081e+17, 1.310674186688705e+17, 1.31067418672933e+17, 1.310674186771517e+17, 1.310674186812142e+17, 1.310674186852768e+17, 1.310674186894956e+17, 1.31067418693558e+17, 1.310674186976205e+17, 1.310674187018392e+17, 1.310674187059018e+17, 1.31067418709808e+17, 1.310674187140268e+17, 1.310674187180892e+17, 1.31067418722933e+17, 1.310674187269955e+17, 1.310674187310579e+17, 1.310674187351205e+17, 1.31067418739183e+17, 1.310674187432454e+17, 1.310674187471517e+17, 1.310674187512142e+17, 1.310674187552767e+17, 1.310674187593393e+17, 1.310674187634017e+17, 1.310674187679331e+17, 1.310674187719955e+17, 1.31067418776058e+17, 1.310674187801204e+17, 1.31067418784183e+17, 1.310674187882455e+17, 1.31067418792308e+17, 1.310674187963706e+17, 1.310674188004329e+17, 1.310674188044955e+17, 1.310674188084018e+17, 1.310674188126204e+17, 1.31067418816683e+17, 1.310674188207455e+17, 1.310674188248081e+17, 1.310674188288705e+17, 1.31067418832933e+17, 1.310674188369956e+17, 1.310674188410579e+17, 1.310674188451205e+17, 1.310674188491831e+17, 1.310674188532454e+17, 1.31067418857308e+17, 1.310674188613705e+17, 1.31067418865433e+17, 1.310674188701204e+17, 1.310674188743392e+17, 1.310674188785581e+17, 1.310674188826205e+17, 1.31067418886683e+17, 1.310674188907455e+17, 1.310674188948081e+17, 1.310674188987142e+17, 1.310674189030892e+17, 1.310674189071517e+17, 1.31067418911058e+17, 1.310674189152767e+17, 1.310674189193393e+17, 1.310674189232456e+17, 1.310674189276205e+17, 1.310674189316829e+17, 1.310674189357455e+17, 1.310674189401204e+17, 1.310674189446518e+17, 1.310674189487142e+17, 1.310674189532454e+17, 1.310674189576205e+17, 1.310674189619955e+17, 1.31067418966058e+17, 1.310674189701204e+17, 1.310674189743393e+17, 1.310674189794956e+17, 1.310674189838705e+17, 1.310674189879331e+17, 1.310674189919955e+17, 1.31067418996058e+17, 1.310674190001204e+17, 1.31067419004183e+17, 1.310674190082455e+17, 1.31067419012308e+17, 1.310674190165267e+17, 1.310674190207455e+17, 1.310674190248081e+17, 1.31067419029183e+17, 1.310674190337142e+17, 1.310674190380893e+17, 1.31067419042308e+17, 1.310674190465267e+17, 1.31067419051058e+17, 1.310674190551205e+17, 1.31067419059183e+17, 1.310674190634017e+17, 1.310674190674643e+17, 1.310674190715268e+17, 1.31067419076058e+17, 1.310674190801204e+17, 1.310674190843393e+17, 1.310674190885581e+17, 1.31067419092933e+17, 1.310674190971517e+17, 1.310674191013705e+17, 1.310674191055892e+17, 1.310674191102767e+17, 1.310674191143392e+17, 1.310674191184018e+17, 1.31067419122933e+17, 1.310674191269955e+17, 1.310674191313705e+17, 1.310674191357455e+17, 1.310674191401206e+17, 1.31067419144183e+17, 1.310674191484017e+17, 1.310674191527767e+17, 1.310674191568393e+17, 1.310674191612142e+17, 1.31067419165433e+17, 1.310674191699643e+17, 1.310674191740268e+17, 1.310674191782455e+17, 1.310674191827768e+17, 1.310674191868392e+17, 1.310674191913705e+17, 1.310674191957455e+17, 1.31067419199808e+17, 1.310674192040268e+17, 1.310674192080892e+17, 1.310674192121517e+17, 1.310674192165267e+17, 1.310674192209018e+17, 1.310674192251205e+17, 1.31067419229183e+17, 1.310674192335579e+17, 1.310674192377768e+17, 1.310674192418392e+17, 1.310674192457454e+17, 1.31067419249808e+17, 1.31067419254183e+17, 1.310674192590267e+17, 1.310674192630893e+17, 1.310674192671517e+17, 1.310674192715268e+17, 1.310674192755892e+17, 1.310674192799643e+17, 1.310674192843392e+17, 1.310674192884018e+17, 1.310674192927767e+17, 1.310674192969956e+17, 1.310674193010579e+17, 1.310674193051205e+17, 1.310674193096517e+17, 1.31067419314183e+17, 1.310674193184018e+17, 1.310674193224643e+17, 1.31067419326683e+17, 1.310674193307455e+17, 1.310674193348081e+17, 1.310674193387142e+17, 1.310674193427767e+17, 1.310674193468393e+17, 1.310674193513705e+17, 1.310674193555892e+17, 1.310674193596517e+17, 1.310674193637143e+17, 1.310674193677768e+17, 1.310674193718392e+17, 1.310674193762143e+17, 1.310674193802767e+17, 1.310674193843393e+17, 1.310674193882455e+17, 1.310674193924643e+17, 1.310674193965268e+17, 1.310674194007455e+17, 1.310674194048079e+17, 1.310674194094956e+17, 1.310674194137143e+17, 1.310674194177768e+17, 1.310674194218392e+17, 1.310674194259017e+17, 1.310674194299643e+17, 1.310674194340268e+17, 1.310674194380892e+17, 1.310674194421518e+17, 1.310674194462141e+17, 1.310674194502767e+17, 1.310674194551205e+17, 1.310674194590267e+17, 1.310674194634017e+17, 1.310674194674642e+17, 1.310674194715268e+17, 1.310674194755892e+17, 1.310674194801204e+17, 1.310674194846518e+17, 1.31067419489183e+17, 1.310674194930893e+17, 1.310674194971517e+17, 1.310674195015268e+17, 1.310674195059018e+17, 1.310674195099642e+17, 1.310674195140268e+17, 1.310674195182455e+17, 1.310674195226204e+17, 1.310674195269955e+17, 1.310674195313705e+17, 1.310674195355892e+17, 1.310674195396517e+17, 1.310674195437143e+17, 1.310674195477768e+17, 1.310674195518392e+17, 1.310674195557455e+17, 1.31067419559808e+17, 1.310674195638705e+17, 1.310674195680892e+17, 1.310674195721518e+17, 1.310674195762143e+17, 1.310674195804329e+17, 1.310674195849642e+17, 1.310674195888704e+17, 1.310674195934017e+17, 1.310674195974642e+17, 1.310674196019955e+17, 1.31067419606058e+17, 1.310674196101204e+17, 1.310674196143392e+17, 1.310674196184018e+17, 1.310674196226205e+17, 1.31067419626683e+17, 1.310674196307455e+17, 1.310674196348081e+17, 1.310674196388705e+17, 1.31067419642933e+17, 1.310674196471517e+17, 1.310674196512143e+17, 1.310674196552768e+17, 1.310674196594954e+17, 1.31067419663558e+17, 1.310674196676205e+17, 1.310674196716831e+17, 1.310674196757454e+17, 1.31067419679808e+17, 1.310674196838706e+17, 1.310674196879329e+17, 1.310674196921517e+17, 1.310674196962143e+17, 1.310674197002767e+17, 1.310674197043392e+17, 1.310674197084017e+17, 1.310674197124643e+17, 1.310674197168393e+17, 1.310674197209018e+17, 1.310674197249642e+17, 1.310674197296517e+17, 1.310674197337143e+17, 1.310674197377766e+17, 1.310674197418392e+17, 1.310674197459018e+17, 1.310674197501206e+17, 1.310674197546516e+17, 1.310674197588705e+17, 1.310674197629331e+17, 1.310674197669955e+17, 1.310674197713705e+17, 1.310674197755892e+17, 1.31067419779808e+17, 1.310674197844955e+17, 1.31067419788558e+17, 1.310674197926205e+17, 1.31067419796683e+17, 1.310674198007455e+17, 1.310674198048081e+17, 1.310674198088704e+17, 1.31067419812933e+17, 1.310674198169956e+17, 1.310674198210579e+17, 1.310674198251205e+17, 1.310674198293393e+17, 1.310674198334017e+17, 1.310674198374642e+17, 1.310674198416829e+17, 1.310674198457455e+17, 1.310674198496517e+17, 1.310674198537143e+17, 1.310674198584018e+17, 1.310674198624643e+17, 1.310674198665267e+17, 1.31067419870433e+17, 1.310674198748081e+17, 1.31067419879183e+17, 1.310674198832456e+17, 1.310674198874643e+17, 1.310674198915268e+17, 1.310674198955892e+17, 1.31067419899808e+17, 1.310674199038706e+17, 1.310674199080893e+17, 1.310674199123081e+17, 1.310674199163704e+17, 1.310674199202769e+17, 1.310674199243392e+17, 1.310674199288705e+17, 1.310674199330893e+17, 1.310674199374642e+17, 1.310674199416831e+17, 1.310674199457455e+17, 1.310674199499643e+17, 1.310674199544955e+17, 1.310674199585581e+17, 1.310674199626204e+17, 1.310674199669956e+17, 1.310674199712143e+17, 1.310674199751205e+17, 1.310674199793393e+17, 1.310674199834019e+17, 1.310674199874642e+17, 1.310674199915268e+17, 1.310674199955892e+17, 1.310674199994954e+17, 1.310674200040268e+17, 1.310674200080892e+17, 1.310674200121518e+17, 1.310674200162143e+17, 1.310674200201204e+17, 1.310674200246518e+17, 1.31067420029183e+17, 1.310674200334017e+17, 1.310674200374643e+17, 1.310674200416831e+17, 1.310674200459018e+17, 1.310674200499643e+17, 1.310674200540268e+17, 1.310674200587142e+17, 1.310674200627767e+17, 1.310674200668393e+17, 1.310674200712142e+17, 1.310674200751205e+17, 1.310674200794956e+17, 1.310674200837143e+17, 1.310674200877768e+17, 1.310674200921518e+17, 1.310674200963706e+17, 1.310674201005893e+17, 1.310674201051205e+17, 1.310674201091831e+17, 1.310674201132454e+17, 1.31067420117308e+17, 1.310674201213705e+17, 1.31067420125433e+17, 1.310674201294956e+17, 1.31067420133558e+17, 1.310674201376205e+17, 1.310674201418392e+17, 1.310674201459017e+17, 1.310674201501204e+17, 1.31067420154183e+17, 1.310674201582455e+17, 1.310674201624643e+17, 1.310674201665267e+17, 1.31067420171058e+17, 1.310674201751205e+17, 1.31067420179183e+17, 1.310674201837142e+17, 1.310674201879329e+17, 1.31067420192308e+17, 1.31067420196683e+17, 1.310674202007455e+17, 1.310674202048079e+17, 1.310674202088705e+17, 1.31067420212933e+17, 1.310674202169955e+17, 1.310674202209018e+17, 1.310674202251205e+17, 1.310674202293393e+17, 1.310674202334017e+17, 1.310674202374643e+17, 1.310674202418392e+17, 1.310674202459017e+17, 1.310674202499642e+17, 1.310674202543393e+17, 1.310674202588704e+17, 1.310674202630893e+17, 1.310674202674642e+17, 1.310674202718392e+17, 1.31067420276058e+17, 1.310674202802767e+17, 1.310674202843392e+17, 1.310674202884018e+17, 1.310674202924643e+17, 1.310674202965267e+17, 1.310674203005893e+17, 1.310674203046518e+17, 1.310674203093393e+17, 1.310674203134017e+17, 1.310674203174643e+17, 1.310674203216829e+17, 1.310674203257455e+17, 1.310674203296518e+17, 1.310674203340268e+17, 1.310674203380892e+17, 1.31067420342308e+17, 1.310674203465267e+17, 1.310674203507455e+17, 1.310674203551205e+17, 1.31067420359183e+17, 1.310674203634017e+17, 1.310674203676205e+17, 1.310674203719955e+17, 1.310674203762143e+17, 1.310674203802767e+17, 1.310674203843393e+17, 1.310674203890267e+17, 1.310674203930893e+17, 1.310674203971517e+17, 1.310674204015268e+17, 1.310674204055892e+17, 1.310674204094956e+17, 1.31067420413558e+17, 1.310674204179331e+17, 1.310674204221518e+17, 1.310674204268393e+17, 1.31067420431058e+17, 1.310674204352767e+17, 1.310674204393393e+17, 1.310674204434017e+17, 1.310674204474643e+17, 1.310674204516829e+17, 1.310674204557454e+17, 1.310674204602767e+17, 1.310674204649642e+17, 1.310674204690268e+17, 1.310674204730893e+17, 1.310674204771517e+17, 1.310674204812142e+17, 1.310674204857455e+17, 1.31067420489808e+17, 1.310674204938705e+17, 1.310674204980892e+17, 1.310674205021518e+17, 1.310674205062143e+17, 1.310674205102767e+17, 1.310674205146518e+17, 1.310674205188704e+17, 1.310674205232454e+17, 1.310674205276205e+17, 1.310674205316829e+17, 1.310674205362143e+17, 1.310674205401204e+17, 1.31067420544183e+17, 1.310674205490268e+17, 1.310674205530893e+17, 1.310674205569956e+17, 1.31067420561058e+17, 1.310674205651204e+17, 1.310674205696517e+17, 1.310674205738706e+17, 1.310674205779329e+17, 1.310674205819955e+17, 1.31067420586058e+17, 1.310674205902769e+17, 1.310674205949642e+17, 1.310674205990267e+17, 1.310674206030893e+17, 1.310674206071517e+17, 1.310674206112142e+17, 1.310674206152768e+17, 1.310674206199643e+17, 1.310674206238705e+17, 1.310674206285581e+17, 1.310674206324643e+17, 1.310674206365268e+17, 1.310674206405892e+17, 1.310674206446516e+17, 1.310674206487142e+17, 1.310674206530893e+17, 1.31067420657308e+17, 1.310674206615268e+17, 1.310674206662143e+17, 1.31067420670433e+17, 1.310674206746518e+17, 1.310674206788705e+17, 1.31067420682933e+17, 1.310674206869955e+17, 1.31067420691058e+17, 1.310674206951205e+17, 1.310674206993393e+17, 1.310674207034017e+17, 1.310674207076205e+17, 1.310674207115268e+17, 1.310674207157455e+17, 1.310674207207455e+17, 1.310674207248079e+17, 1.310674207293393e+17, 1.310674207334017e+17, 1.310674207376205e+17, 1.310674207418392e+17, 1.310674207459018e+17, 1.310674207499643e+17, 1.310674207541829e+17, 1.310674207582455e+17, 1.310674207624643e+17, 1.31067420766683e+17, 1.310674207707456e+17, 1.310674207748079e+17, 1.310674207788704e+17, 1.31067420782933e+17, 1.310674207869955e+17, 1.310674207912142e+17, 1.310674207951205e+17, 1.310674207993393e+17, 1.31067420803558e+17, 1.310674208074643e+17, 1.310674208116829e+17, 1.310674208157455e+17, 1.310674208196517e+17, 1.310674208237143e+17, 1.310674208279331e+17, 1.31067420832308e+17, 1.310674208363706e+17, 1.310674208405893e+17, 1.310674208446516e+17, 1.310674208487142e+17, 1.31067420852933e+17, 1.31067420857308e+17, 1.310674208619955e+17, 1.31067420866058e+17, 1.310674208702767e+17, 1.310674208744955e+17, 1.310674208788705e+17, 1.31067420882933e+17, 1.310674208869956e+17, 1.31067420891058e+17, 1.310674208951205e+17, 1.31067420899183e+17, 1.310674209032456e+17, 1.31067420907308e+17, 1.310674209113705e+17, 1.31067420915433e+17, 1.310674209196518e+17, 1.310674209237142e+17, 1.310674209277768e+17, 1.310674209318392e+17, 1.310674209360581e+17, 1.310674209401204e+17, 1.310674209441829e+17, 1.310674209484018e+17, 1.310674209524643e+17, 1.31067420956683e+17, 1.310674209609018e+17, 1.310674209649642e+17, 1.310674209690267e+17, 1.310674209732456e+17, 1.31067420977308e+17, 1.310674209813705e+17, 1.31067420985433e+17, 1.310674209896517e+17, 1.310674209937143e+17, 1.310674209977766e+17, 1.310674210016831e+17, 1.310674210059018e+17, 1.310674210099642e+17, 1.310674210140268e+17, 1.310674210180892e+17, 1.310674210219955e+17, 1.31067421026058e+17, 1.310674210301206e+17, 1.31067421034183e+17, 1.310674210382455e+17, 1.310674210423081e+17, 1.310674210462143e+17, 1.310674210509018e+17, 1.310674210549642e+17, 1.310674210590267e+17, 1.310674210640268e+17, 1.310674210682455e+17, 1.31067421072933e+17, 1.310674210769956e+17, 1.31067421081058e+17, 1.310674210852767e+17, 1.310674210893393e+17, 1.31067421093558e+17, 1.310674210977768e+17, 1.310674211019955e+17, 1.31067421106058e+17, 1.310674211099643e+17, 1.310674211143392e+17, 1.310674211184017e+17, 1.310674211224643e+17, 1.310674211263704e+17, 1.310674211305893e+17, 1.310674211346518e+17, 1.310674211387142e+17, 1.31067421142933e+17, 1.310674211469956e+17, 1.31067421151058e+17, 1.310674211552768e+17, 1.310674211593393e+17, 1.310674211634017e+17, 1.310674211674643e+17, 1.310674211715267e+17, 1.310674211762143e+17, 1.31067421180433e+17, 1.310674211851205e+17, 1.310674211894956e+17, 1.310674211937143e+17, 1.310674211977768e+17, 1.310674212018392e+17, 1.310674212059017e+17, 1.310674212102767e+17, 1.310674212143392e+17, 1.310674212184018e+17, 1.31067421222933e+17, 1.310674212269956e+17, 1.310674212313705e+17, 1.310674212355892e+17, 1.310674212402767e+17, 1.310674212444955e+17, 1.310674212487142e+17, 1.310674212527767e+17, 1.310674212571516e+17, 1.310674212612142e+17, 1.310674212652768e+17, 1.31067421269183e+17, 1.310674212732456e+17, 1.310674212774643e+17, 1.310674212815268e+17, 1.310674212857455e+17, 1.31067421289808e+17, 1.310674212937143e+17, 1.310674212977768e+17, 1.310674213023081e+17, 1.310674213062143e+17, 1.310674213105892e+17, 1.310674213146518e+17, 1.310674213188705e+17, 1.31067421322933e+17, 1.31067421327308e+17, 1.310674213318392e+17, 1.310674213362143e+17, 1.310674213402767e+17, 1.310674213443393e+17, 1.310674213484018e+17, 1.310674213524643e+17, 1.31067421356683e+17, 1.310674213607456e+17, 1.310674213648081e+17, 1.310674213693393e+17, 1.31067421373558e+17, 1.310674213776206e+17, 1.310674213816829e+17, 1.31067421386058e+17, 1.310674213901204e+17, 1.31067421394183e+17, 1.310674213984018e+17, 1.310674214027767e+17, 1.310674214068393e+17, 1.310674214109018e+17, 1.310674214154331e+17, 1.310674214194956e+17, 1.31067421423558e+17, 1.310674214277768e+17, 1.310674214318392e+17, 1.310674214357455e+17, 1.310674214402769e+17, 1.310674214443392e+17, 1.31067421448558e+17, 1.310674214526205e+17, 1.31067421456683e+17, 1.310674214612142e+17, 1.31067421465433e+17, 1.310674214694956e+17, 1.310674214737143e+17, 1.310674214777768e+17, 1.310674214818392e+17, 1.31067421486058e+17, 1.310674214901204e+17, 1.310674214946516e+17, 1.310674214988705e+17, 1.31067421502933e+17, 1.31067421507308e+17, 1.310674215113705e+17, 1.310674215152768e+17, 1.310674215194954e+17, 1.310674215234017e+17, 1.310674215276205e+17, 1.310674215316829e+17, 1.310674215357455e+17, 1.310674215402767e+17, 1.31067421544183e+17, 1.310674215490268e+17, 1.310674215534017e+17, 1.310674215577768e+17, 1.310674215619955e+17, 1.31067421566058e+17, 1.310674215701204e+17, 1.310674215744956e+17, 1.31067421578558e+17, 1.310674215830893e+17, 1.310674215871517e+17, 1.310674215913705e+17, 1.31067421595433e+17, 1.310674215996517e+17, 1.310674216037143e+17, 1.310674216079331e+17, 1.31067421612308e+17, 1.310674216168392e+17, 1.310674216209018e+17, 1.310674216251205e+17, 1.310674216294954e+17, 1.31067421633558e+17, 1.310674216376206e+17, 1.310674216418392e+17, 1.310674216459017e+17, 1.310674216499643e+17, 1.310674216540268e+17, 1.310674216580892e+17, 1.310674216619955e+17, 1.310674216662143e+17, 1.310674216701204e+17, 1.31067421674183e+17, 1.310674216784018e+17, 1.31067421682308e+17, 1.310674216863704e+17, 1.31067421690433e+17, 1.310674216944955e+17, 1.310674216987142e+17, 1.310674217027767e+17, 1.310674217068393e+17, 1.310674217113705e+17, 1.310674217154331e+17, 1.310674217194954e+17, 1.310674217237142e+17, 1.310674217277768e+17, 1.310674217318394e+17, 1.310674217359017e+17, 1.31067421739808e+17, 1.310674217444955e+17, 1.310674217488705e+17, 1.31067421753558e+17, 1.310674217576205e+17, 1.310674217616831e+17, 1.310674217659017e+17, 1.310674217699643e+17, 1.310674217741829e+17, 1.310674217785581e+17, 1.310674217826204e+17, 1.310674217865268e+17, 1.31067421791058e+17, 1.310674217951205e+17, 1.31067421799183e+17, 1.31067421803558e+17, 1.310674218077768e+17, 1.310674218119955e+17, 1.31067421816058e+17, 1.310674218202767e+17, 1.310674218243393e+17, 1.310674218284018e+17, 1.310674218324643e+17, 1.31067421840433e+17, 1.310674218444955e+17, 1.310674218487142e+17, 1.31067421852933e+17, 1.310674218569956e+17, 1.310674218610579e+17, 1.310674218651205e+17, 1.31067421869183e+17, 1.310674218734017e+17, 1.310674218774642e+17, 1.310674218815268e+17, 1.310674218855892e+17, 1.310674218896517e+17, 1.310674218937143e+17, 1.310674218977768e+17, 1.310674219018392e+17, 1.310674219057455e+17, 1.310674219099643e+17, 1.310674219146518e+17, 1.310674219187142e+17, 1.310674219226205e+17, 1.31067421926683e+17, 1.310674219307455e+17, 1.310674219348081e+17, 1.310674219387142e+17, 1.31067421942933e+17, 1.310674219469955e+17, 1.310674219513705e+17, 1.310674219555892e+17, 1.310674219596518e+17, 1.310674219637142e+17, 1.310674219677768e+17, 1.310674219719955e+17, 1.310674219768393e+17, 1.310674219813705e+17, 1.31067421985433e+17, 1.310674219894956e+17, 1.31067421993558e+17, 1.310674219979331e+17, 1.310674220019955e+17, 1.310674220062141e+17, 1.31067422010433e+17, 1.310674220144955e+17, 1.310674220187142e+17, 1.310674220227768e+17, 1.31067422026683e+17, 1.310674220307456e+17, 1.310674220348079e+17, 1.310674220388704e+17, 1.31067422042933e+17, 1.310674220469955e+17, 1.310674220516829e+17, 1.310674220559017e+17, 1.31067422060433e+17, 1.310674220644955e+17, 1.310674220684018e+17, 1.310674220727767e+17, 1.31067422076683e+17, 1.310674220807455e+17, 1.310674220849642e+17, 1.310674220890268e+17, 1.310674220930892e+17, 1.31067422097308e+17, 1.310674221015267e+17, 1.310674221054331e+17, 1.310674221096518e+17, 1.310674221137142e+17, 1.310674221177768e+17, 1.310674221218392e+17, 1.310674221257455e+17, 1.31067422130433e+17, 1.310674221348079e+17, 1.310674221388705e+17, 1.310674221432454e+17, 1.31067422147308e+17, 1.310674221519955e+17, 1.31067422156058e+17, 1.310674221601204e+17, 1.310674221641829e+17, 1.310674221682455e+17, 1.310674221723081e+17, 1.31067422176683e+17, 1.310674221807456e+17, 1.310674221848079e+17, 1.310674221890267e+17, 1.310674221930893e+17, 1.310674221971517e+17, 1.310674222012142e+17, 1.31067422206058e+17, 1.310674222101204e+17, 1.31067422214183e+17, 1.310674222184018e+17, 1.310674222224643e+17, 1.31067422226683e+17, 1.310674222313705e+17, 1.310674222354331e+17, 1.310674222394954e+17, 1.310674222434017e+17, 1.310674222482455e+17, 1.31067422252308e+17, 1.310674222563704e+17, 1.31067422260433e+17, 1.310674222649642e+17, 1.310674222693393e+17, 1.310674222737143e+17, 1.310674222779331e+17, 1.310674222819954e+17, 1.31067422286058e+17, 1.310674222905892e+17, 1.310674222946518e+17, 1.310674222987142e+17, 1.310674223027767e+17, 1.310674223074642e+17, 1.310674223115268e+17, 1.310674223159017e+17, 1.310674223201204e+17, 1.310674223249642e+17, 1.310674223290268e+17, 1.310674223330893e+17, 1.310674223371517e+17, 1.310674223412142e+17, 1.310674223452767e+17, 1.310674223493393e+17, 1.310674223534017e+17, 1.31067422357308e+17, 1.310674223615267e+17, 1.310674223659017e+17, 1.310674223702769e+17, 1.310674223746518e+17, 1.310674223788705e+17, 1.310674223830893e+17, 1.310674223871517e+17, 1.310674223912142e+17, 1.31067422395433e+17, 1.310674223994956e+17, 1.310674224037143e+17, 1.310674224079331e+17, 1.310674224121518e+17, 1.31067422416683e+17, 1.310674224209018e+17, 1.310674224249644e+17, 1.310674224290267e+17, 1.310674224330893e+17, 1.31067422437308e+17, 1.310674224412142e+17, 1.310674224452768e+17, 1.310674224501204e+17, 1.310674224540268e+17, 1.310674224580892e+17, 1.310674224626205e+17, 1.310674224665267e+17, 1.310674224709016e+17, 1.310674224754331e+17, 1.310674224794954e+17, 1.31067422483558e+17, 1.310674224876205e+17, 1.310674224916829e+17, 1.310674224957455e+17, 1.31067422500433e+17, 1.310674225049642e+17, 1.310674225090268e+17, 1.310674225130893e+17, 1.310674225177768e+17, 1.310674225218392e+17, 1.310674225259018e+17, 1.310674225302767e+17, 1.310674225343393e+17, 1.310674225387142e+17, 1.310674225430893e+17, 1.31067422547308e+17, 1.310674225513705e+17, 1.31067422555433e+17, 1.310674225596517e+17, 1.310674225638705e+17, 1.310674225679331e+17, 1.310674225719955e+17, 1.31067422576058e+17, 1.310674225801204e+17, 1.310674225848081e+17, 1.310674225890268e+17, 1.310674225934017e+17, 1.310674225977768e+17, 1.310674226018392e+17, 1.310674226059017e+17, 1.310674226101204e+17, 1.310674226143392e+17, 1.310674226184018e+17, 1.310674226224643e+17, 1.310674226265267e+17, 1.310674226307455e+17, 1.310674226348081e+17, 1.310674226387142e+17, 1.310674226427767e+17, 1.310674226469955e+17, 1.31067422651058e+17, 1.310674226549642e+17, 1.31067422659183e+17, 1.310674226630893e+17, 1.310674226679331e+17, 1.310674226727768e+17, 1.310674226768392e+17, 1.310674226809018e+17, 1.310674226849644e+17, 1.310674226893393e+17, 1.310674226934017e+17, 1.310674226974642e+17, 1.310674227016829e+17, 1.310674227057455e+17, 1.310674227096517e+17, 1.310674227138705e+17, 1.310674227179331e+17, 1.310674227226205e+17, 1.310674227265267e+17, 1.310674227305893e+17, 1.310674227348081e+17, 1.310674227388704e+17, 1.31067422742933e+17, 1.310674227469956e+17, 1.310674227510579e+17, 1.310674227551205e+17, 1.31067422759183e+17, 1.310674227630892e+17, 1.310674227671517e+17, 1.310674227712143e+17, 1.310674227752768e+17, 1.31067422779808e+17, 1.310674227848081e+17, 1.310674227890268e+17, 1.310674227934017e+17, 1.310674227974643e+17, 1.310674228018392e+17, 1.310674228059017e+17, 1.310674228099642e+17, 1.310674228143393e+17, 1.310674228184017e+17, 1.310674228227767e+17, 1.310674228269955e+17, 1.310674228312142e+17, 1.310674228355892e+17, 1.310674228396517e+17, 1.31067422844183e+17, 1.310674228482455e+17, 1.310674228526205e+17, 1.31067422856683e+17, 1.310674228609018e+17, 1.310674228649642e+17, 1.310674228690268e+17, 1.310674228730892e+17, 1.310674228769956e+17, 1.310674228821517e+17, 1.310674228863704e+17, 1.31067422890433e+17, 1.310674228944955e+17, 1.31067422898558e+17, 1.310674229026205e+17, 1.31067422906683e+17, 1.310674229107455e+17, 1.310674229149642e+17, 1.310674229190268e+17, 1.310674229232456e+17, 1.31067422927308e+17, 1.310674229313705e+17, 1.310674229355892e+17, 1.31067422939808e+17, 1.310674229441829e+17, 1.31067422948558e+17, 1.310674229530893e+17, 1.310674229571517e+17, 1.310674229612142e+17, 1.31067422965433e+17, 1.310674229694956e+17, 1.31067422973558e+17, 1.310674229776205e+17, 1.310674229816831e+17, 1.310674229855892e+17, 1.310674229899643e+17, 1.310674229940268e+17, 1.310674229980892e+17, 1.310674230021518e+17, 1.310674230068392e+17, 1.310674230109018e+17, 1.310674230148081e+17, 1.31067423019183e+17, 1.310674230232454e+17, 1.31067423027308e+17, 1.310674230316829e+17, 1.310674230359017e+17, 1.310674230399643e+17, 1.310674230443392e+17, 1.31067423048558e+17, 1.310674230565267e+17, 1.310674230609018e+17, 1.310674230651205e+17, 1.31067423069183e+17, 1.310674230734017e+17, 1.310674230774643e+17, 1.310674230815268e+17, 1.310674230859018e+17, 1.310674230899643e+17, 1.310674230940268e+17, 1.310674230980893e+17, 1.310674231023081e+17, 1.310674231063704e+17, 1.31067423110433e+17, 1.310674231143392e+17, 1.310674231187142e+17, 1.310674231226205e+17, 1.31067423126683e+17, 1.310674231309018e+17, 1.310674231349642e+17, 1.310674231390268e+17, 1.31067423142933e+17, 1.310674231469955e+17, 1.31067423151058e+17, 1.310674231551205e+17, 1.31067423159183e+17, 1.310674231632456e+17, 1.31067423167308e+17, 1.310674231713705e+17, 1.31067423175433e+17, 1.31067423179808e+17, 1.310674231838705e+17, 1.310674231887142e+17, 1.310674231927767e+17, 1.310674231968392e+17, 1.310674232009018e+17, 1.310674232049642e+17, 1.310674232088705e+17, 1.310674232129331e+17, 1.310674232169955e+17, 1.310674232213705e+17, 1.31067423225433e+17, 1.310674232294956e+17, 1.310674232338705e+17, 1.310674232379331e+17, 1.310674232419955e+17, 1.310674232465267e+17, 1.310674232510579e+17, 1.310674232555892e+17, 1.31067423259808e+17, 1.31067423264183e+17, 1.310674232690267e+17, 1.310674232730893e+17, 1.31067423277308e+17, 1.310674232816831e+17, 1.310674232859017e+17, 1.310674232901206e+17, 1.310674232943393e+17, 1.310674232988704e+17, 1.31067423302933e+17, 1.310674233069955e+17, 1.31067423311058e+17, 1.310674233152767e+17, 1.310674233191831e+17, 1.31067423324183e+17, 1.310674233282455e+17, 1.31067423332308e+17, 1.310674233363706e+17, 1.31067423340433e+17, 1.310674233444955e+17, 1.31067423348558e+17, 1.310674233526205e+17, 1.31067423356683e+17, 1.310674233607455e+17, 1.310674233646518e+17, 1.310674233690268e+17, 1.310674233730893e+17, 1.310674233773079e+17, 1.310674233813705e+17, 1.310674233857455e+17, 1.31067423389808e+17, 1.310674233938705e+17, 1.310674233980892e+17, 1.31067423402308e+17, 1.31067423406683e+17, 1.310674234107455e+17, 1.310674234148081e+17, 1.310674234188705e+17, 1.31067423422933e+17, 1.310674234274643e+17, 1.310674234315268e+17, 1.310674234355892e+17, 1.310674234396517e+17, 1.310674234437143e+17, 1.310674234477768e+17, 1.310674234518392e+17, 1.310674234559018e+17, 1.310674234601206e+17, 1.310674234641829e+17, 1.310674234682455e+17, 1.310674234723081e+17, 1.310674234763704e+17, 1.31067423480433e+17, 1.310674234844955e+17, 1.310674234884017e+17, 1.310674234924643e+17, 1.310674234965267e+17, 1.310674235007455e+17, 1.310674235048079e+17, 1.310674235088705e+17, 1.31067423512933e+17, 1.310674235169955e+17, 1.31067423521058e+17, 1.310674235252768e+17, 1.310674235293393e+17, 1.310674235334017e+17, 1.310674235376205e+17, 1.310674235416831e+17, 1.310674235457455e+17, 1.310674235501206e+17, 1.310674235541829e+17, 1.310674235582455e+17, 1.31067423562308e+17, 1.310674235663704e+17, 1.31067423570433e+17, 1.310674235744955e+17, 1.310674235788705e+17, 1.310674235829331e+17, 1.310674235869955e+17, 1.310674235910579e+17, 1.31067423596058e+17, 1.310674236001204e+17, 1.310674236044955e+17, 1.31067423608558e+17, 1.310674236130892e+17, 1.310674236176205e+17, 1.310674236216831e+17, 1.310674236257455e+17, 1.310674236299642e+17, 1.310674236338705e+17, 1.310674236380892e+17, 1.310674236426205e+17, 1.31067423646683e+17, 1.310674236509018e+17, 1.310674236549642e+17, 1.31067423659183e+17, 1.310674236634017e+17, 1.310674236679331e+17, 1.310674236721518e+17, 1.310674236762141e+17, 1.310674236802767e+17, 1.310674236843393e+17, 1.310674236888705e+17, 1.310674236927768e+17, 1.310674236968393e+17, 1.310674237009018e+17, 1.31067423705433e+17, 1.310674237094954e+17, 1.31067423713558e+17, 1.310674237174642e+17, 1.310674237218392e+17, 1.310674237262143e+17, 1.31067423730433e+17, 1.310674237344955e+17, 1.310674237385581e+17, 1.310674237427767e+17, 1.310674237471517e+17, 1.310674237515268e+17, 1.310674237557454e+17, 1.310674237599643e+17, 1.310674237640268e+17, 1.310674237680892e+17, 1.310674237721517e+17, 1.310674237762143e+17, 1.310674237802767e+17, 1.31067423784183e+17, 1.31067423788558e+17, 1.310674237926205e+17, 1.31067423796683e+17, 1.31067423801058e+17, 1.310674238051205e+17, 1.31067423809183e+17, 1.310674238134017e+17, 1.310674238174643e+17, 1.310674238219955e+17, 1.310674238265268e+17, 1.310674238305892e+17, 1.310674238352767e+17, 1.310674238393393e+17, 1.310674238434017e+17, 1.310674238474642e+17, 1.310674238518392e+17, 1.310674238557455e+17, 1.31067423860433e+17, 1.310674238644955e+17, 1.31067423868558e+17, 1.310674238726205e+17, 1.310674238765267e+17, 1.31067423881058e+17, 1.310674238851205e+17, 1.310674238894954e+17, 1.31067423893558e+17, 1.310674238976205e+17, 1.310674239016829e+17, 1.310674239062143e+17, 1.310674239109018e+17, 1.310674239149642e+17, 1.310674239190268e+17, 1.310674239230893e+17, 1.31067423927308e+17, 1.310674239315268e+17, 1.310674239355892e+17, 1.310674239396517e+17, 1.310674239435579e+17, 1.310674239477768e+17, 1.310674239518392e+17, 1.310674239559017e+17, 1.310674239601206e+17, 1.31067423964183e+17, 1.310674239684017e+17, 1.310674239724643e+17, 1.310674239765268e+17, 1.310674239807455e+17, 1.310674239848079e+17, 1.310674239888705e+17, 1.310674239930893e+17, 1.310674239971517e+17, 1.310674240013705e+17, 1.31067424005433e+17, 1.310674240096517e+17, 1.310674240137143e+17, 1.310674240176205e+17, 1.310674240216831e+17, 1.31067424026058e+17, 1.310674240301206e+17, 1.31067424034183e+17, 1.310674240387142e+17, 1.310674240432454e+17, 1.310674240476206e+17, 1.310674240516829e+17, 1.310674240557455e+17, 1.310674240596517e+17, 1.310674240638705e+17, 1.310674240679331e+17, 1.31067424072308e+17, 1.310674240763706e+17, 1.31067424080433e+17, 1.310674240849642e+17, 1.31067424089183e+17, 1.310674240932456e+17, 1.310674240974643e+17, 1.310674241015267e+17, 1.31067424105433e+17, 1.310674241096518e+17, 1.31067424113558e+17, 1.310674241176205e+17, 1.310674241216831e+17, 1.310674241257454e+17, 1.310674241302767e+17, 1.310674241343392e+17, 1.310674241384018e+17, 1.310674241426204e+17, 1.310674241465267e+17, 1.310674241505892e+17, 1.310674241546518e+17, 1.310674241596517e+17, 1.310674241637143e+17, 1.310674241679331e+17, 1.310674241721518e+17, 1.310674241765267e+17, 1.310674241805893e+17, 1.310674241846518e+17, 1.310674241885581e+17, 1.310674241926204e+17, 1.31067424196683e+17, 1.310674242009018e+17, 1.310674242052767e+17, 1.310674242099643e+17, 1.310674242140268e+17, 1.310674242179331e+17, 1.310674242224643e+17, 1.310674242265267e+17, 1.31067424230433e+17, 1.310674242344955e+17, 1.31067424238558e+17, 1.310674242427768e+17, 1.310674242468393e+17, 1.310674242513705e+17, 1.310674242557455e+17, 1.310674242601204e+17, 1.310674242643392e+17, 1.310674242687142e+17, 1.310674242727767e+17, 1.310674242768393e+17, 1.31067424281058e+17, 1.310674242851205e+17, 1.31067424289183e+17, 1.31067424293558e+17, 1.310674242976205e+17, 1.31067424302308e+17, 1.310674243063706e+17, 1.31067424310433e+17, 1.310674243149644e+17, 1.310674243190267e+17, 1.31067424322933e+17, 1.310674243271517e+17, 1.310674243312142e+17, 1.310674243352768e+17, 1.31067424339183e+17, 1.310674243432454e+17, 1.310674243476205e+17, 1.31067424352308e+17, 1.310674243563704e+17, 1.31067424361058e+17, 1.310674243651205e+17, 1.310674243694956e+17, 1.310674243738705e+17, 1.310674243779329e+17, 1.310674243819955e+17, 1.310674243862143e+17, 1.310674243902767e+17, 1.310674243946518e+17, 1.310674243987142e+17, 1.310674244034017e+17, 1.310674244076205e+17, 1.310674244116829e+17, 1.31067424416058e+17, 1.310674244201204e+17, 1.31067424424183e+17, 1.310674244282455e+17, 1.310674244323081e+17, 1.310674244365267e+17, 1.310674244409018e+17, 1.310674244449642e+17, 1.310674244490267e+17, 1.310674244530893e+17, 1.310674244574642e+17, 1.310674244616829e+17, 1.31067424466058e+17, 1.310674244701204e+17, 1.310674244743392e+17, 1.310674244784018e+17, 1.310674244824643e+17, 1.310674244866829e+17, 1.310674244907455e+17, 1.310674244949642e+17, 1.310674244990268e+17, 1.310674245030892e+17, 1.310674245071517e+17, 1.310674245112143e+17, 1.310674245154331e+17, 1.310674245194954e+17, 1.31067424523558e+17, 1.310674245287142e+17, 1.310674245327767e+17, 1.310674245368393e+17, 1.310674245409018e+17, 1.310674245455892e+17, 1.310674245496517e+17, 1.310674245538705e+17, 1.310674245580893e+17, 1.310674245624643e+17, 1.310674245665268e+17, 1.310674245705893e+17, 1.310674245744955e+17, 1.310674245785581e+17, 1.310674245832454e+17, 1.31067424587308e+17, 1.310674245913705e+17, 1.31067424595433e+17, 1.310674245994954e+17, 1.31067424603558e+17, 1.310674246077768e+17, 1.310674246118392e+17, 1.310674246159017e+17, 1.310674246199643e+17, 1.310674246238705e+17, 1.310674246279331e+17, 1.31067424632308e+17, 1.310674246363706e+17, 1.310674246407455e+17, 1.310674246448081e+17, 1.310674246493393e+17, 1.310674246534017e+17, 1.310674246574642e+17, 1.310674246616829e+17, 1.310674246659017e+17, 1.310674246701204e+17, 1.310674246744955e+17, 1.31067424678558e+17, 1.310674246832456e+17, 1.310674246874643e+17, 1.310674246915268e+17, 1.310674246955892e+17, 1.310674246996517e+17, 1.310674247037143e+17, 1.310674247079331e+17, 1.310674247119955e+17, 1.310674247159018e+17, 1.310674247201206e+17, 1.310674247241829e+17, 1.310674247282455e+17, 1.310674247324643e+17, 1.310674247365268e+17, 1.310674247405892e+17, 1.310674247448079e+17, 1.310674247488705e+17, 1.31067424752933e+17, 1.310674247569955e+17, 1.310674247613705e+17, 1.310674247657455e+17, 1.31067424769808e+17, 1.310674247740268e+17, 1.310674247787142e+17, 1.310674247830893e+17, 1.310674247871517e+17, 1.310674247912143e+17, 1.310674247954331e+17, 1.310674247999643e+17, 1.310674248040268e+17, 1.310674248080892e+17, 1.310674248121517e+17, 1.310674248162143e+17, 1.310674248202767e+17, 1.310674248243392e+17, 1.310674248284018e+17, 1.310674248326205e+17, 1.310674248369955e+17, 1.310674248412143e+17, 1.31067424845433e+17, 1.310674248494956e+17, 1.31067424853558e+17, 1.310674248576205e+17, 1.310674248616831e+17, 1.310674248657454e+17, 1.310674248701206e+17, 1.310674248741829e+17, 1.310674248787142e+17, 1.310674248827767e+17, 1.310674248871517e+17, 1.310674248915268e+17, 1.310674248957455e+17, 1.31067424899808e+17, 1.310674249038705e+17, 1.310674249080892e+17, 1.310674249121518e+17, 1.310674249163706e+17, 1.310674249204329e+17, 1.310674249248081e+17, 1.310674249288704e+17, 1.31067424932933e+17, 1.31067424937308e+17, 1.310674249413705e+17, 1.31067424945433e+17, 1.310674249499643e+17, 1.310674249540269e+17, 1.310674249582455e+17, 1.31067424962308e+17, 1.310674249663706e+17, 1.31067424970433e+17, 1.310674249746518e+17, 1.310674249788705e+17, 1.310674249827768e+17, 1.310674249869955e+17, 1.310674249915267e+17, 1.310674249955892e+17, 1.310674249996518e+17, 1.310674250037142e+17, 1.310674250079329e+17, 1.310674250119955e+17, 1.310674250160581e+17, 1.310674250199643e+17, 1.310674250240268e+17, 1.310674250282455e+17, 1.310674250321517e+17, 1.310674250362143e+17, 1.310674250402769e+17, 1.310674250443392e+17, 1.310674250487142e+17, 1.310674250527767e+17, 1.310674250568393e+17, 1.310674250612142e+17, 1.310674250652768e+17, 1.310674250693393e+17, 1.310674250734017e+17, 1.310674250777766e+17, 1.310674250819955e+17, 1.31067425086058e+17, 1.310674250907455e+17, 1.310674250949644e+17, 1.310674250991831e+17, 1.310674251034017e+17, 1.310674251076205e+17, 1.310674251116829e+17, 1.31067425116058e+17, 1.310674251201204e+17, 1.31067425124183e+17, 1.310674251287142e+17, 1.31067425132933e+17, 1.310674251369955e+17, 1.31067425141058e+17, 1.310674251451205e+17, 1.31067425149183e+17, 1.310674251534017e+17, 1.310674251576205e+17, 1.310674251619955e+17, 1.31067425166683e+17, 1.310674251707455e+17, 1.310674251751205e+17, 1.31067425179183e+17, 1.310674251832454e+17, 1.310674251871517e+17, 1.310674251913705e+17, 1.31067425195433e+17, 1.310674251993393e+17, 1.31067425203558e+17, 1.310674252082455e+17, 1.310674252127768e+17, 1.310674252171517e+17, 1.310674252212142e+17, 1.31067425225433e+17, 1.310674252294954e+17, 1.31067425233558e+17, 1.310674252379331e+17, 1.310674252421518e+17, 1.310674252463704e+17, 1.31067425250433e+17, 1.310674252544955e+17, 1.310674252585581e+17, 1.310674252626205e+17, 1.31067425266683e+17, 1.310674252707455e+17, 1.310674252748081e+17, 1.310674252788704e+17, 1.310674252827768e+17, 1.310674252869956e+17, 1.310674252912143e+17, 1.310674252952767e+17, 1.31067425299808e+17, 1.310674253038705e+17, 1.310674253079329e+17, 1.310674253119955e+17, 1.31067425316058e+17, 1.310674253199643e+17, 1.310674253243392e+17, 1.310674253284018e+17, 1.310674253326205e+17, 1.310674253369955e+17, 1.31067425341058e+17, 1.310674253451205e+17, 1.31067425349183e+17, 1.310674253532456e+17, 1.31067425357308e+17, 1.310674253618392e+17, 1.310674253659018e+17, 1.310674253699642e+17, 1.310674253743392e+17, 1.310674253787144e+17, 1.310674253830893e+17, 1.310674253871517e+17, 1.310674253912142e+17, 1.310674253952768e+17, 1.310674253993393e+17, 1.310674254032454e+17, 1.310674254074643e+17, 1.310674254118392e+17, 1.310674254159017e+17, 1.310674254199643e+17, 1.310674254244955e+17, 1.310674254285581e+17, 1.310674254326205e+17, 1.31067425437308e+17, 1.310674254418394e+17, 1.310674254463704e+17, 1.310674254507455e+17, 1.310674254548081e+17, 1.310674254588705e+17, 1.310674254630893e+17, 1.310674254671517e+17, 1.310674254712143e+17, 1.310674254752768e+17, 1.310674254805892e+17, 1.310674254848079e+17, 1.310674254893393e+17, 1.310674254934017e+17, 1.310674254974642e+17, 1.310674255015268e+17, 1.31067425505433e+17, 1.310674255094956e+17, 1.310674255146518e+17, 1.310674255187142e+17, 1.310674255227767e+17, 1.310674255268393e+17, 1.310674255309018e+17, 1.310674255349642e+17, 1.310674255390268e+17, 1.310674255430892e+17, 1.310674255471517e+17, 1.310674255510579e+17, 1.310674255551205e+17, 1.310674255596518e+17, 1.310674255640268e+17, 1.310674255680892e+17, 1.310674255726205e+17, 1.310674255768393e+17, 1.310674255809018e+17, 1.310674255857455e+17, 1.310674255901206e+17, 1.310674255941829e+17, 1.310674255984017e+17, 1.310674256024643e+17, 1.310674256065268e+17, 1.310674256105892e+17, 1.310674256146516e+17, 1.31067425618558e+17, 1.310674256226204e+17, 1.310674256269955e+17, 1.310674256312142e+17, 1.310674256352768e+17, 1.310674256396517e+17, 1.310674256437143e+17, 1.310674256477768e+17, 1.310674256521518e+17, 1.310674256565267e+17, 1.310674256605893e+17, 1.310674256685581e+17, 1.310674256726205e+17, 1.31067425676683e+17, 1.310674256807455e+17, 1.310674256849644e+17, 1.310674256888705e+17, 1.310674256932454e+17, 1.31067425697308e+17, 1.310674257016829e+17, 1.310674257059017e+17, 1.310674257101204e+17, 1.31067425714183e+17, 1.310674257184018e+17, 1.310674257226205e+17, 1.31067425726683e+17, 1.310674257307455e+17, 1.310674257349642e+17, 1.310674257390268e+17, 1.31067425742933e+17, 1.310674257469956e+17, 1.31067425751058e+17, 1.310674257551204e+17, 1.31067425759183e+17, 1.310674257632456e+17, 1.310674257674643e+17, 1.310674257715267e+17, 1.310674257755892e+17, 1.310674257796518e+17, 1.310674257837142e+17, 1.310674257879329e+17, 1.310674257919955e+17, 1.310674257959017e+17, 1.310674257999643e+17, 1.310674258040268e+17, 1.310674258084018e+17, 1.310674258124643e+17, 1.310674258165267e+17, 1.310674258213705e+17, 1.31067425825433e+17, 1.310674258294956e+17, 1.31067425833558e+17, 1.310674258382455e+17, 1.310674258423081e+17, 1.310674258465267e+17, 1.310674258505892e+17, 1.310674258546518e+17, 1.310674258591831e+17, 1.310674258632454e+17, 1.310674258679329e+17, 1.310674258719955e+17, 1.31067425876058e+17, 1.310674258801204e+17, 1.31067425884183e+17, 1.310674258882455e+17, 1.310674258924643e+17, 1.31067425896683e+17, 1.310674259015268e+17, 1.310674259060581e+17, 1.310674259101204e+17, 1.310674259141829e+17, 1.310674259182455e+17, 1.310674259224643e+17, 1.310674259268393e+17, 1.310674259315268e+17, 1.310674259357455e+17, 1.31067425939808e+17, 1.310674259438705e+17, 1.310674259482455e+17, 1.310674259523081e+17, 1.310674259565267e+17, 1.310674259605893e+17, 1.310674259644955e+17, 1.310674259687142e+17, 1.310674259727768e+17, 1.31067425976683e+17, 1.310674259809018e+17, 1.310674259849644e+17, 1.310674259890267e+17, 1.310674259934017e+17, 1.310674259974642e+17, 1.310674260015268e+17, 1.310674260059017e+17, 1.310674260101204e+17, 1.310674260148081e+17, 1.310674260190268e+17, 1.31067426022933e+17, 1.310674260274643e+17, 1.310674260315267e+17, 1.310674260355892e+17, 1.310674260401204e+17, 1.31067426044183e+17, 1.310674260490267e+17, 1.310674260530893e+17, 1.31067426057308e+17, 1.310674260618392e+17, 1.310674260659017e+17, 1.310674260699643e+17, 1.310674260743393e+17, 1.310674260784018e+17, 1.310674260824643e+17, 1.310674260863706e+17, 1.31067426090433e+17, 1.310674260948079e+17, 1.310674260990267e+17, 1.310674261030893e+17, 1.310674261071517e+17, 1.310674261112142e+17, 1.310674261152768e+17, 1.310674261194954e+17, 1.31067426123558e+17, 1.310674261280892e+17, 1.310674261324643e+17, 1.31067426136683e+17, 1.310674261412143e+17, 1.310674261452768e+17, 1.310674261493393e+17, 1.31067426153558e+17, 1.310674261576205e+17, 1.310674261618392e+17, 1.310674261659017e+17, 1.310674261699643e+17, 1.310674261738706e+17, 1.310674261782455e+17, 1.31067426182308e+17, 1.310674261863704e+17, 1.31067426190433e+17, 1.310674261944955e+17, 1.310674261988705e+17, 1.31067426202933e+17, 1.310674262069955e+17, 1.310674262112142e+17, 1.310674262155892e+17, 1.310674262196517e+17, 1.310674262238705e+17, 1.310674262279331e+17, 1.310674262321518e+17, 1.31067426236683e+17, 1.310674262407455e+17, 1.310674262449644e+17, 1.310674262488705e+17, 1.310674262534017e+17, 1.310674262577768e+17, 1.310674262621517e+17, 1.310674262663706e+17, 1.31067426270433e+17, 1.310674262744955e+17, 1.310674262784018e+17, 1.310674262824643e+17, 1.310674262865267e+17, 1.310674262905893e+17, 1.310674262948081e+17, 1.310674262988704e+17, 1.31067426302933e+17, 1.310674263069956e+17, 1.310674263110579e+17, 1.310674263155892e+17, 1.310674263196517e+17, 1.310674263238705e+17, 1.310674263279331e+17, 1.310674263324643e+17, 1.310674263369955e+17, 1.31067426341058e+17, 1.310674263451205e+17, 1.31067426349183e+17, 1.310674263532456e+17, 1.31067426357308e+17, 1.310674263619954e+17, 1.31067426366058e+17, 1.310674263701206e+17, 1.31067426374183e+17, 1.310674263784017e+17, 1.310674263824643e+17, 1.310674263865268e+17, 1.310674263909018e+17, 1.310674263949642e+17, 1.310674263996517e+17, 1.310674264037143e+17, 1.310674264080892e+17, 1.310674264124643e+17, 1.310674264171517e+17, 1.310674264212143e+17, 1.310674264252767e+17, 1.310674264293393e+17, 1.310674264334017e+17, 1.310674264376205e+17, 1.310674264416829e+17, 1.310674264459017e+17, 1.310674264499643e+17, 1.31067426454183e+17, 1.310674264584017e+17, 1.310674264624643e+17, 1.310674264665267e+17, 1.310674264705893e+17, 1.310674264746518e+17, 1.310674264787142e+17, 1.31067426486683e+17, 1.310674264907455e+17, 1.310674264948081e+17, 1.310674264988705e+17, 1.310674265032456e+17, 1.31067426507308e+17, 1.310674265112143e+17, 1.31067426515433e+17, 1.310674265194956e+17, 1.31067426523558e+17, 1.310674265276205e+17, 1.310674265321517e+17, 1.310674265360581e+17, 1.310674265402767e+17, 1.310674265443392e+17, 1.310674265484018e+17, 1.310674265524643e+17, 1.310674265565267e+17, 1.310674265607455e+17, 1.310674265648081e+17, 1.310674265688705e+17, 1.31067426572933e+17, 1.310674265769955e+17, 1.310674265812142e+17, 1.310674265852768e+17, 1.310674265893393e+17, 1.310674265934017e+17, 1.31067426597308e+17, 1.310674266016831e+17, 1.310674266059018e+17, 1.31067426610433e+17, 1.310674266146516e+17, 1.310674266190267e+17, 1.310674266230893e+17, 1.310674266271517e+17, 1.310674266319955e+17, 1.310674266365267e+17, 1.310674266409018e+17, 1.310674266452768e+17, 1.310674266493393e+17, 1.310674266543392e+17, 1.310674266584017e+17, 1.310674266624643e+17, 1.310674266669955e+17, 1.310674266709018e+17, 1.31067426675433e+17, 1.310674266799643e+17, 1.310674266840268e+17, 1.310674266880892e+17, 1.310674266921518e+17, 1.310674266962143e+17, 1.310674267002767e+17, 1.310674267046516e+17, 1.310674267087142e+17, 1.310674267127768e+17, 1.31067426716683e+17, 1.310674267209018e+17, 1.310674267249644e+17, 1.31067426729183e+17, 1.310674267332454e+17, 1.310674267376205e+17, 1.310674267415268e+17, 1.310674267496517e+17, 1.310674267537143e+17, 1.310674267577768e+17, 1.310674267618392e+17, 1.31067426766058e+17, 1.310674267702767e+17, 1.310674267744955e+17, 1.310674267787142e+17, 1.310674267827767e+17, 1.310674267868393e+17, 1.31067426791058e+17, 1.310674267951204e+17, 1.31067426799183e+17, 1.310674268030892e+17, 1.310674268071517e+17, 1.310674268112143e+17, 1.310674268152767e+17, 1.310674268194954e+17, 1.31067426823558e+17, 1.310674268276205e+17, 1.31067426832308e+17, 1.31067426836683e+17, 1.310674268409018e+17, 1.310674268451205e+17, 1.310674268493393e+17, 1.310674268534017e+17, 1.310674268582455e+17, 1.310674268626204e+17, 1.31067426866683e+17, 1.310674268707455e+17, 1.310674268746516e+17, 1.310674268787142e+17, 1.310674268827767e+17, 1.310674268869955e+17, 1.310674268910579e+17, 1.310674268951205e+17, 1.31067426899183e+17, 1.310674269034017e+17, 1.310674269074642e+17, 1.310674269115268e+17, 1.310674269155892e+17, 1.310674269196517e+17, 1.31067426923558e+17, 1.310674269276205e+17, 1.310674269316829e+17, 1.31067426936683e+17, 1.310674269407455e+17, 1.310674269446516e+17, 1.310674269487142e+17, 1.310674269530892e+17, 1.310674269571517e+17, 1.310674269613705e+17, 1.310674269657455e+17, 1.310674269701204e+17, 1.310674269746518e+17, 1.310674269787142e+17, 1.310674269827767e+17, 1.310674269868393e+17, 1.310674269909018e+17, 1.310674269949642e+17, 1.310674269988705e+17, 1.31067427002933e+17, 1.310674270069956e+17, 1.31067427011058e+17, 1.310674270152768e+17, 1.310674270193393e+17, 1.310674270234017e+17, 1.310674270274643e+17, 1.310674270315267e+17, 1.310674270355892e+17, 1.310674270399642e+17, 1.310674270440268e+17, 1.310674270480893e+17, 1.310674270521517e+17, 1.310674270562143e+17, 1.310674270605892e+17, 1.310674270646518e+17, 1.310674270687142e+17, 1.310674270730893e+17, 1.310674270771517e+17, 1.310674270812142e+17, 1.310674270852768e+17, 1.310674270893393e+17, 1.310674270934017e+17, 1.310674270974642e+17, 1.310674271015268e+17, 1.310674271059017e+17, 1.31067427109808e+17, 1.310674271138705e+17, 1.310674271179331e+17, 1.310674271219955e+17, 1.31067427126058e+17, 1.310674271301204e+17, 1.310674271341829e+17, 1.310674271380892e+17, 1.310674271421517e+17, 1.310674271462143e+17, 1.31067427150433e+17, 1.310674271544955e+17, 1.310674271587144e+17, 1.310674271627767e+17, 1.310674271668392e+17, 1.310674271709018e+17, 1.310674271749642e+17, 1.310674271790267e+17, 1.310674271830893e+17, 1.310674271871517e+17, 1.310674271912142e+17, 1.31067427196058e+17, 1.310674272001204e+17, 1.310674272040268e+17, 1.310674272085581e+17, 1.310674272126205e+17, 1.31067427216683e+17, 1.310674272205893e+17, 1.310674272248081e+17, 1.310674272288704e+17, 1.31067427232933e+17, 1.310674272369956e+17, 1.310674272413705e+17, 1.31067427245433e+17, 1.310674272496517e+17, 1.31067427254183e+17, 1.310674272582455e+17, 1.31067427262933e+17, 1.310674272669956e+17, 1.310674272712142e+17, 1.310674272754331e+17, 1.31067427279808e+17, 1.310674272840268e+17, 1.310674272882455e+17, 1.310674272926204e+17, 1.31067427296683e+17, 1.310674273007455e+17, 1.310674273046518e+17, 1.310674273090267e+17, 1.310674273130893e+17, 1.310674273171517e+17, 1.310674273212142e+17, 1.310674273252768e+17, 1.310674273293393e+17, 1.310674273334017e+17, 1.310674273376205e+17, 1.310674273416829e+17, 1.310674273457455e+17, 1.310674273496517e+17, 1.310674273544955e+17, 1.310674273587142e+17, 1.310674273627768e+17, 1.310674273669956e+17, 1.310674273713705e+17, 1.31067427375433e+17, 1.310674273796517e+17, 1.310674273837143e+17, 1.31067427388558e+17, 1.310674273926205e+17, 1.310674273965267e+17, 1.310674274005893e+17, 1.310674274046518e+17, 1.310674274088705e+17, 1.31067427412933e+17, 1.310674274169956e+17, 1.31067427421058e+17, 1.310674274252768e+17, 1.310674274293393e+17, 1.310674274334017e+17, 1.310674274377768e+17, 1.310674274416831e+17, 1.310674274459017e+17, 1.310674274499642e+17, 1.310674274540268e+17, 1.310674274580892e+17, 1.310674274624643e+17, 1.31067427466683e+17, 1.310674274705893e+17, 1.310674274746518e+17, 1.310674274790268e+17, 1.310674274830893e+17, 1.310674274871517e+17, 1.310674274916831e+17, 1.310674274959018e+17, 1.310674274999643e+17, 1.310674275041829e+17, 1.310674275087142e+17, 1.310674275127768e+17, 1.310674275168393e+17, 1.310674275215268e+17, 1.310674275262143e+17, 1.310674275302767e+17, 1.310674275344955e+17, 1.310674275390268e+17, 1.310674275430893e+17, 1.310674275480893e+17, 1.310674275521517e+17, 1.310674275562143e+17, 1.310674275607455e+17, 1.310674275648079e+17, 1.310674275690267e+17, 1.310674275730893e+17, 1.310674275771517e+17, 1.310674275813705e+17, 1.310674275859017e+17, 1.310674275902767e+17, 1.310674275943393e+17, 1.310674275984018e+17, 1.310674276024643e+17, 1.310674276065268e+17, 1.310674276107455e+17, 1.310674276149644e+17, 1.310674276190267e+17, 1.310674276230893e+17, 1.31067427627308e+17, 1.310674276313705e+17, 1.31067427635433e+17, 1.310674276396517e+17, 1.310674276437143e+17, 1.310674276477768e+17, 1.310674276521518e+17, 1.310674276562143e+17, 1.310674276602767e+17, 1.310674276643392e+17, 1.310674276685581e+17, 1.310674276726205e+17, 1.31067427676683e+17, 1.310674276807455e+17, 1.310674276848081e+17, 1.310674276888704e+17, 1.31067427692933e+17, 1.310674276971517e+17, 1.310674277012143e+17, 1.310674277052767e+17, 1.310674277093393e+17, 1.310674277134017e+17, 1.310674277174642e+17, 1.310674277226205e+17, 1.310674277268393e+17, 1.31067427731058e+17, 1.310674277355892e+17, 1.31067427739808e+17, 1.310674277443393e+17, 1.310674277484017e+17, 1.310674277527768e+17, 1.310674277568392e+17, 1.310674277609018e+17, 1.31067427765433e+17, 1.310674277694956e+17, 1.310674277737142e+17, 1.310674277777768e+17, 1.310674277819955e+17, 1.310674277865267e+17, 1.310674277909018e+17, 1.310674277949642e+17, 1.310674277993393e+17, 1.310674278034017e+17, 1.310674278076205e+17, 1.310674278116831e+17, 1.310674278157455e+17, 1.310674278202769e+17, 1.310674278243392e+17, 1.310674278284017e+17, 1.310674278326205e+17, 1.310674278368393e+17, 1.310674278409018e+17, 1.310674278455892e+17, 1.310674278496517e+17, 1.310674278538705e+17, 1.310674278579331e+17, 1.310674278619955e+17, 1.310674278662141e+17, 1.310674278702767e+17, 1.310674278744955e+17, 1.310674278785581e+17, 1.310674278827768e+17, 1.310674278868393e+17, 1.310674278910579e+17, 1.31067427895433e+17, 1.310674278996517e+17, 1.310674279037143e+17, 1.310674279077768e+17, 1.310674279119955e+17, 1.31067427916058e+17, 1.310674279201204e+17, 1.310674279240268e+17, 1.310674279284018e+17, 1.310674279324643e+17, 1.310674279363706e+17, 1.31067427940433e+17, 1.310674279451204e+17, 1.31067427949183e+17, 1.310674279532456e+17, 1.310674279576205e+17, 1.310674279616829e+17, 1.310674279655892e+17, 1.310674279699643e+17, 1.310674279740268e+17, 1.310674279782455e+17, 1.310674279824643e+17, 1.310674279868393e+17, 1.310674279912142e+17, 1.31067427995433e+17, 1.310674279994956e+17, 1.310674280038705e+17, 1.310674280080893e+17, 1.310674280121518e+17, 1.310674280162143e+17, 1.31067428020433e+17, 1.310674280243393e+17, 1.310674280285581e+17, 1.310674280326204e+17, 1.310674280371517e+17, 1.310674280412142e+17, 1.31067428045433e+17, 1.310674280496517e+17, 1.310674280537143e+17, 1.310674280577768e+17, 1.310674280619955e+17, 1.310674280663704e+17, 1.310674280707455e+17, 1.310674280748081e+17, 1.310674280788704e+17, 1.310674280834017e+17, 1.310674280874643e+17, 1.310674280915268e+17, 1.310674280962143e+17, 1.310674281001204e+17, 1.310674281046518e+17, 1.310674281088705e+17, 1.310674281130893e+17, 1.310674281171517e+17, 1.310674281215268e+17, 1.310674281257455e+17, 1.31067428129808e+17, 1.310674281340268e+17, 1.310674281380892e+17, 1.310674281421518e+17, 1.310674281463706e+17, 1.31067428150433e+17, 1.310674281544955e+17, 1.310674281585581e+17, 1.310674281632454e+17, 1.31067428167308e+17, 1.310674281716829e+17, 1.310674281759017e+17, 1.310674281799643e+17, 1.310674281840268e+17, 1.310674281880892e+17, 1.310674281921517e+17, 1.310674281962143e+17, 1.31067428200433e+17, 1.310674282044955e+17, 1.310674282093393e+17, 1.31067428213558e+17, 1.310674282180892e+17, 1.310674282219955e+17, 1.310674282262143e+17, 1.310674282309018e+17, 1.310674282349642e+17, 1.310674282390267e+17, 1.310674282430893e+17, 1.310674282471517e+17, 1.310674282512142e+17, 1.310674282551205e+17, 1.31067428259183e+17, 1.31067428263558e+17, 1.310674282677766e+17, 1.310674282718392e+17, 1.310674282759018e+17, 1.310674282802767e+17, 1.310674282843393e+17, 1.310674282885581e+17, 1.310674282926204e+17, 1.310674282968393e+17, 1.310674283013705e+17, 1.31067428305433e+17, 1.310674283094956e+17, 1.310674283137143e+17, 1.310674283179331e+17, 1.310674283221518e+17, 1.310674283262143e+17, 1.310674283302767e+17, 1.310674283382455e+17, 1.31067428342933e+17, 1.310674283469956e+17, 1.310674283510579e+17, 1.310674283551205e+17, 1.31067428359183e+17, 1.310674283632454e+17, 1.310674283676205e+17, 1.310674283716829e+17, 1.310674283757455e+17, 1.310674283799643e+17, 1.31067428384183e+17, 1.310674283882455e+17, 1.31067428392308e+17, 1.310674283971517e+17, 1.310674284019955e+17, 1.310674284063704e+17, 1.31067428410433e+17, 1.310674284144955e+17, 1.310674284185581e+17, 1.310674284226204e+17, 1.31067428426683e+17, 1.310674284307456e+17, 1.310674284349642e+17, 1.310674284390267e+17, 1.310674284430893e+17, 1.310674284476205e+17, 1.310674284518392e+17, 1.31067428456058e+17, 1.310674284601204e+17, 1.310674284648081e+17, 1.310674284693393e+17, 1.310674284734017e+17, 1.310674284774642e+17, 1.310674284821517e+17, 1.310674284862143e+17, 1.310674284902767e+17, 1.310674284946518e+17, 1.310674284990267e+17, 1.310674285032456e+17, 1.31067428507308e+17, 1.310674285113704e+17, 1.310674285155892e+17, 1.310674285196517e+17, 1.310674285237143e+17, 1.310674285282455e+17, 1.31067428532308e+17, 1.310674285363704e+17, 1.31067428540433e+17, 1.310674285444955e+17, 1.310674285484017e+17, 1.310674285526204e+17, 1.31067428556683e+17, 1.310674285613705e+17, 1.31067428565433e+17, 1.310674285694956e+17, 1.31067428573558e+17, 1.310674285776205e+17, 1.310674285816831e+17, 1.310674285857455e+17, 1.31067428589808e+17, 1.310674285938705e+17, 1.310674285979331e+17, 1.310674286018392e+17, 1.310674286062143e+17, 1.310674286102767e+17, 1.310674286143393e+17, 1.310674286190268e+17, 1.310674286232454e+17, 1.31067428627308e+17, 1.310674286315268e+17, 1.310674286359017e+17, 1.310674286402767e+17, 1.310674286443392e+17, 1.310674286484018e+17, 1.310674286524643e+17, 1.310674286565267e+17, 1.310674286605893e+17, 1.310674286649642e+17, 1.310674286690268e+17, 1.310674286730893e+17, 1.31067428677308e+17, 1.310674286813705e+17, 1.310674286854331e+17, 1.310674286894956e+17, 1.31067428693558e+17, 1.310674286980893e+17, 1.310674287021517e+17, 1.310674287065267e+17, 1.310674287109018e+17, 1.310674287149642e+17, 1.310674287193393e+17, 1.31067428723558e+17, 1.310674287277768e+17, 1.310674287321518e+17, 1.310674287362143e+17, 1.310674287402767e+17, 1.310674287443393e+17, 1.310674287484018e+17, 1.310674287524643e+17, 1.310674287568392e+17, 1.310674287610579e+17, 1.31067428765433e+17, 1.310674287693393e+17, 1.310674287734019e+17, 1.310674287779331e+17, 1.310674287819955e+17, 1.310674287862143e+17, 1.310674287907455e+17, 1.310674287948081e+17, 1.310674287990268e+17, 1.310674288032456e+17, 1.310674288076205e+17, 1.310674288116831e+17, 1.310674288157455e+17, 1.310674288201206e+17, 1.310674288248079e+17, 1.310674288288705e+17, 1.31067428832933e+17, 1.31067428837308e+17, 1.310674288413705e+17, 1.31067428845433e+17, 1.310674288494956e+17, 1.31067428854183e+17, 1.310674288587142e+17, 1.31067428862933e+17, 1.310674288669956e+17, 1.310674288713705e+17, 1.310674288754331e+17, 1.310674288794956e+17, 1.310674288837142e+17, 1.310674288877768e+17, 1.310674288918392e+17, 1.310674288959017e+17, 1.31067428899808e+17, 1.310674289038705e+17, 1.310674289080892e+17, 1.310674289121518e+17, 1.310674289162143e+17, 1.310674289202767e+17, 1.310674289243392e+17, 1.310674289285581e+17, 1.310674289324643e+17, 1.31067428936683e+17, 1.310674289409018e+17, 1.310674289449642e+17, 1.310674289490268e+17, 1.310674289532456e+17, 1.310674289576205e+17, 1.310674289619955e+17, 1.310674289662143e+17, 1.310674289702769e+17, 1.310674289743392e+17, 1.310674289784017e+17, 1.310674289826205e+17, 1.310674289868393e+17, 1.310674289909018e+17, 1.310674289952768e+17, 1.310674289993393e+17, 1.310674290034017e+17, 1.310674290074643e+17, 1.310674290116831e+17, 1.310674290157455e+17, 1.31067429019808e+17, 1.310674290237143e+17, 1.310674290279331e+17, 1.310674290318392e+17, 1.310674290359017e+17, 1.310674290399642e+17, 1.310674290440268e+17, 1.310674290480893e+17, 1.310674290524643e+17, 1.310674290565268e+17, 1.310674290605892e+17, 1.310674290646516e+17, 1.310674290687142e+17, 1.310674290727767e+17, 1.310674290768393e+17, 1.310674290809018e+17, 1.310674290852768e+17, 1.310674290893393e+17, 1.310674290934017e+17, 1.310674290980892e+17, 1.310674291021518e+17, 1.310674291062143e+17, 1.310674291101206e+17, 1.31067429114183e+17, 1.310674291182455e+17, 1.31067429122308e+17, 1.310674291265268e+17, 1.310674291307455e+17, 1.310674291348081e+17, 1.310674291388705e+17, 1.310674291432454e+17, 1.310674291471517e+17, 1.310674291516829e+17, 1.310674291562143e+17, 1.310674291607455e+17, 1.310674291648081e+17, 1.310674291688705e+17, 1.31067429172933e+17, 1.310674291769955e+17, 1.31067429181058e+17, 1.310674291852768e+17, 1.310674291894956e+17, 1.31067429193558e+17, 1.310674291976205e+17, 1.310674292016831e+17, 1.310674292057454e+17, 1.31067429209808e+17, 1.310674292137142e+17, 1.310674292177768e+17, 1.310674292221517e+17, 1.310674292262143e+17, 1.310674292302769e+17, 1.310674292343392e+17, 1.310674292384017e+17, 1.310674292424643e+17, 1.31067429246683e+17, 1.310674292507455e+17, 1.310674292548079e+17, 1.310674292587142e+17, 1.310674292627767e+17, 1.31067429267308e+17, 1.310674292713705e+17, 1.31067429275433e+17, 1.31067429279808e+17, 1.310674292837143e+17, 1.310674292880892e+17, 1.310674292921518e+17, 1.310674292963704e+17, 1.31067429300433e+17, 1.310674293044955e+17, 1.310674293085581e+17, 1.310674293127767e+17, 1.310674293169955e+17, 1.310674293212142e+17, 1.310674293255892e+17, 1.310674293296517e+17, 1.310674293337143e+17, 1.310674293380892e+17, 1.310674293424643e+17, 1.310674293469956e+17, 1.31067429351058e+17, 1.310674293555892e+17, 1.310674293596517e+17, 1.310674293640268e+17, 1.310674293684018e+17, 1.310674293724643e+17, 1.310674293765267e+17, 1.310674293809018e+17, 1.310674293849642e+17, 1.310674293890267e+17, 1.310674293932456e+17, 1.31067429397308e+17, 1.310674294013704e+17, 1.31067429405433e+17, 1.310674294094956e+17, 1.31067429413558e+17, 1.310674294176205e+17, 1.310674294216831e+17, 1.310674294265268e+17, 1.310674294309018e+17, 1.310674294352767e+17, 1.310674294393393e+17, 1.310674294434017e+17, 1.310674294474642e+17, 1.310674294519955e+17, 1.310674294565267e+17, 1.310674294609018e+17, 1.310674294648081e+17, 1.310674294688705e+17, 1.31067429472933e+17, 1.310674294769955e+17, 1.31067429481058e+17, 1.310674294851205e+17, 1.310674294894954e+17, 1.310674294938705e+17, 1.310674294980892e+17, 1.31067429502308e+17, 1.310674295065267e+17, 1.310674295107455e+17, 1.310674295157455e+17, 1.310674295199643e+17, 1.310674295240268e+17, 1.310674295285581e+17, 1.31067429532933e+17, 1.310674295369956e+17, 1.310674295416829e+17, 1.310674295457455e+17, 1.310674295502767e+17, 1.310674295544955e+17, 1.310674295590268e+17, 1.310674295634017e+17, 1.310674295674643e+17, 1.310674295715268e+17, 1.310674295755892e+17, 1.310674295796517e+17, 1.310674295837142e+17, 1.310674295877768e+17, 1.310674295916831e+17, 1.310674295963704e+17, 1.31067429600433e+17, 1.310674296043392e+17, 1.31067429608558e+17, 1.310674296124643e+17, 1.31067429616683e+17, 1.310674296207455e+17, 1.310674296248079e+17, 1.310674296288705e+17, 1.310674296327767e+17, 1.310674296368393e+17, 1.310674296409018e+17, 1.310674296449642e+17, 1.310674296490267e+17, 1.310674296530893e+17, 1.310674296571517e+17, 1.310674296612142e+17, 1.310674296655892e+17, 1.310674296696517e+17, 1.310674296737143e+17, 1.310674296779331e+17, 1.310674296819955e+17, 1.310674296859018e+17, 1.310674296899643e+17, 1.310674296941829e+17, 1.310674296982455e+17, 1.310674297027767e+17, 1.310674297068393e+17, 1.310674297110579e+17, 1.310674297152768e+17, 1.310674297193393e+17, 1.310674297234017e+17, 1.310674297279331e+17, 1.310674297321518e+17, 1.310674297365267e+17, 1.310674297405893e+17, 1.310674297446516e+17, 1.310674297487142e+17, 1.310674297526205e+17, 1.310674297576205e+17, 1.310674297616829e+17, 1.310674297663704e+17, 1.310674297707455e+17, 1.31067429775433e+17, 1.310674297794956e+17, 1.310674297834017e+17, 1.310674297874643e+17, 1.310674297916831e+17, 1.31067429796058e+17, 1.310674298001204e+17, 1.310674298049644e+17, 1.310674298091831e+17, 1.31067429813558e+17, 1.310674298177768e+17, 1.310674298218392e+17, 1.310674298259017e+17, 1.310674298299643e+17, 1.310674298340268e+17, 1.310674298380892e+17, 1.31067429842308e+17, 1.310674298463704e+17, 1.31067429850433e+17, 1.310674298544955e+17, 1.310674298587142e+17, 1.310674298627767e+17, 1.310674298668393e+17, 1.310674298712143e+17, 1.310674298752767e+17, 1.310674298793393e+17, 1.310674298840268e+17, 1.310674298880892e+17, 1.310674298921517e+17, 1.31067429896058e+17, 1.310674299001204e+17, 1.31067429904183e+17, 1.310674299082455e+17, 1.31067429912308e+17, 1.310674299165267e+17, 1.310674299205893e+17, 1.310674299244955e+17, 1.310674299290268e+17, 1.310674299332456e+17, 1.31067429937308e+17, 1.310674299415268e+17, 1.310674299457454e+17, 1.31067429949808e+17, 1.310674299548079e+17, 1.310674299588705e+17, 1.310674299630893e+17, 1.31067429967308e+17, 1.310674299713705e+17, 1.310674299755892e+17, 1.310674299796517e+17, 1.310674299837143e+17, 1.310674299879331e+17, 1.310674299919955e+17, 1.31067429996058e+17, 1.310674299999643e+17, 1.31067430004183e+17, 1.310674300082455e+17, 1.31067430012308e+17, 1.310674300162141e+17, 1.310674300205893e+17, 1.310674300246516e+17, 1.310674300290267e+17, 1.310674300340268e+17, 1.31067430038558e+17, 1.310674300426205e+17, 1.310674300469955e+17, 1.310674300513705e+17, 1.310674300559018e+17, 1.310674300599642e+17, 1.310674300640268e+17, 1.310674300680892e+17, 1.310674300721517e+17, 1.310674300763704e+17, 1.310674300805892e+17, 1.310674300852768e+17, 1.310674300896517e+17, 1.310674300937143e+17, 1.310674300977768e+17, 1.310674301019955e+17, 1.310674301062143e+17, 1.310674301102767e+17, 1.310674301144955e+17, 1.310674301185581e+17, 1.310674301226205e+17, 1.310674301269956e+17, 1.310674301316829e+17, 1.310674301359017e+17, 1.31067430139808e+17, 1.310674301443392e+17, 1.310674301488705e+17, 1.31067430152933e+17, 1.310674301571517e+17, 1.310674301615268e+17, 1.310674301655892e+17, 1.31067430169808e+17, 1.310674301737143e+17, 1.310674301782455e+17, 1.310674301823081e+17, 1.310674301865267e+17, 1.310674301905892e+17, 1.310674301946518e+17, 1.310674301987142e+17, 1.310674302027767e+17, 1.310674302068392e+17, 1.310674302109018e+17, 1.310674302149642e+17, 1.310674302190267e+17, 1.310674302229331e+17, 1.310674302269955e+17, 1.310674302312142e+17, 1.31067430236058e+17, 1.310674302401204e+17, 1.31067430244183e+17, 1.31067430248558e+17, 1.31067430252933e+17, 1.31067430257308e+17, 1.310674302612143e+17, 1.310674302654331e+17, 1.31067430269808e+17, 1.310674302738705e+17, 1.310674302779329e+17, 1.310674302821517e+17, 1.310674302862143e+17, 1.310674302902767e+17, 1.310674302946518e+17, 1.310674302987142e+17, 1.310674303027767e+17, 1.310674303069955e+17, 1.31067430311058e+17, 1.310674303149642e+17, 1.310674303193393e+17, 1.310674303234017e+17, 1.310674303274643e+17, 1.310674303318392e+17, 1.310674303359018e+17, 1.310674303401206e+17, 1.310674303443392e+17, 1.310674303484017e+17, 1.310674303526205e+17, 1.31067430356683e+17, 1.310674303612142e+17, 1.31067430365433e+17, 1.310674303694956e+17, 1.310674303738705e+17, 1.310674303779331e+17, 1.310674303819955e+17, 1.31067430386058e+17, 1.310674303901204e+17, 1.31067430394183e+17, 1.310674303984018e+17, 1.310674304024643e+17, 1.310674304063706e+17, 1.310674304104329e+17, 1.310674304146518e+17, 1.310674304185581e+17, 1.310674304226204e+17, 1.31067430427308e+17, 1.310674304318392e+17, 1.310674304357455e+17, 1.31067430439808e+17, 1.31067430444183e+17, 1.310674304488705e+17, 1.310674304530893e+17, 1.31067430457308e+17, 1.310674304615268e+17, 1.310674304659018e+17, 1.310674304699643e+17, 1.310674304740268e+17, 1.310674304780893e+17, 1.310674304821517e+17, 1.310674304863704e+17, 1.310674304909018e+17, 1.310674304952768e+17, 1.310674304994956e+17, 1.31067430503558e+17, 1.310674305077768e+17, 1.310674305118392e+17, 1.310674305159017e+17, 1.310674305199643e+17, 1.310674305240268e+17, 1.310674305280892e+17, 1.310674305321518e+17, 1.310674305362141e+17, 1.310674305405893e+17, 1.310674305448081e+17, 1.310674305488705e+17, 1.310674305527768e+17, 1.310674305574642e+17, 1.310674305615268e+17, 1.310674305659017e+17, 1.310674305699643e+17, 1.31067430574183e+17, 1.310674305784018e+17, 1.310674305826205e+17, 1.31067430586683e+17, 1.310674305909016e+17, 1.310674305952768e+17, 1.310674305994956e+17, 1.31067430603558e+17, 1.310674306076205e+17, 1.310674306118392e+17, 1.310674306159018e+17, 1.310674306199643e+17, 1.310674306246518e+17, 1.310674306287142e+17, 1.310674306332454e+17, 1.31067430637308e+17, 1.310674306415268e+17, 1.310674306459018e+17, 1.310674306499643e+17, 1.31067430654183e+17, 1.310674306584018e+17, 1.31067430662933e+17, 1.310674306671517e+17, 1.310674306712143e+17, 1.310674306752768e+17, 1.31067430679808e+17, 1.310674306838705e+17, 1.310674306879329e+17, 1.310674306921518e+17, 1.310674306962143e+17, 1.310674307002767e+17, 1.310674307048081e+17, 1.310674307088705e+17, 1.31067430712933e+17, 1.310674307169956e+17, 1.31067430721058e+17, 1.310674307259018e+17, 1.310674307302767e+17, 1.310674307343392e+17, 1.310674307384017e+17, 1.310674307426204e+17, 1.31067430746683e+17, 1.310674307507455e+17, 1.310674307548081e+17, 1.310674307593393e+17, 1.310674307634017e+17, 1.310674307674642e+17, 1.310674307716831e+17, 1.310674307757455e+17, 1.31067430779808e+17, 1.310674307838705e+17, 1.310674307879331e+17, 1.310674307919955e+17, 1.31067430796058e+17, 1.310674308001204e+17, 1.310674308043393e+17, 1.310674308084017e+17, 1.310674308124643e+17, 1.31067430816683e+17, 1.310674308207456e+17, 1.310674308252768e+17, 1.310674308294954e+17, 1.31067430833558e+17, 1.310674308379329e+17, 1.310674308421518e+17, 1.310674308463704e+17, 1.310674308509016e+17, 1.310674308551205e+17, 1.31067430859183e+17, 1.310674308632456e+17, 1.310674308673079e+17, 1.310674308712142e+17, 1.310674308754331e+17, 1.310674308793393e+17, 1.310674308834017e+17, 1.310674308874643e+17, 1.310674308915267e+17, 1.31067430896058e+17, 1.310674309002769e+17, 1.310674309043392e+17, 1.310674309088705e+17, 1.310674309127767e+17, 1.310674309168393e+17, 1.310674309213704e+17, 1.31067430925433e+17, 1.310674309294956e+17, 1.31067430933558e+17, 1.310674309376205e+17, 1.310674309418392e+17, 1.310674309459018e+17, 1.310674309501204e+17, 1.310674309541829e+17, 1.310674309584017e+17, 1.310674309630893e+17, 1.310674309669955e+17, 1.310674309710579e+17, 1.310674309751205e+17, 1.31067430979183e+17, 1.310674309834017e+17, 1.310674309876205e+17, 1.310674309916831e+17, 1.310674309962143e+17, 1.31067431000433e+17, 1.310674310044955e+17, 1.310674310090268e+17, 1.31067431013558e+17, 1.310674310176205e+17, 1.310674310219955e+17, 1.310674310260581e+17, 1.310674310305893e+17, 1.310674310349642e+17, 1.310674310390268e+17, 1.310674310430893e+17, 1.310674310471517e+17, 1.31067431051058e+17, 1.310674310551205e+17, 1.31067431059183e+17, 1.310674310632456e+17, 1.310674310679331e+17, 1.310674310719954e+17, 1.31067431076058e+17, 1.310674310801206e+17, 1.310674310844955e+17, 1.310674310885581e+17, 1.310674310930893e+17, 1.310674310971517e+17, 1.310674311015268e+17, 1.310674311059017e+17, 1.310674311099643e+17, 1.310674311140268e+17, 1.310674311180892e+17, 1.310674311224643e+17, 1.31067431126683e+17, 1.310674311307455e+17, 1.310674311348081e+17, 1.310674311388704e+17, 1.31067431142933e+17, 1.310674311469956e+17, 1.310674311510579e+17, 1.310674311551205e+17, 1.310674311594954e+17, 1.31067431163558e+17, 1.310674311679329e+17, 1.310674311719955e+17, 1.31067431176058e+17, 1.310674311799643e+17, 1.31067431184183e+17, 1.310674311880892e+17, 1.310674311927767e+17, 1.310674311968393e+17, 1.310674312009018e+17, 1.310674312052768e+17, 1.310674312094956e+17, 1.310674312138705e+17, 1.310674312179331e+17, 1.310674312219955e+17, 1.310674312265268e+17, 1.310674312309018e+17, 1.310674312352768e+17, 1.310674312394956e+17, 1.31067431243558e+17, 1.310674312476205e+17, 1.310674312516831e+17, 1.310674312557455e+17, 1.31067431259808e+17, 1.310674312638705e+17, 1.310674312679331e+17, 1.31067431272308e+17, 1.310674312765267e+17, 1.310674312805893e+17, 1.310674312849644e+17, 1.310674312890268e+17, 1.310674312932454e+17, 1.31067431297308e+17, 1.310674313013705e+17, 1.31067431305433e+17, 1.31067431309808e+17, 1.310674313144955e+17, 1.310674313187142e+17, 1.310674313226205e+17, 1.310674313268393e+17, 1.310674313309018e+17, 1.310674313349642e+17, 1.310674313390268e+17, 1.310674313432456e+17, 1.31067431347308e+17, 1.310674313516831e+17, 1.310674313557454e+17, 1.31067431359808e+17, 1.310674313638706e+17, 1.310674313679329e+17, 1.310674313719955e+17, 1.31067431376058e+17, 1.310674313802769e+17, 1.310674313843392e+17, 1.310674313884017e+17, 1.310674313924643e+17, 1.31067431396683e+17, 1.310674314007455e+17, 1.310674314048079e+17, 1.31067431409183e+17, 1.310674314132454e+17, 1.310674314179331e+17, 1.310674314221518e+17, 1.31067431426683e+17, 1.310674314310579e+17, 1.310674314351205e+17, 1.31067431439183e+17, 1.310674314434019e+17, 1.310674314474642e+17, 1.310674314515268e+17, 1.31067431456058e+17, 1.310674314601204e+17, 1.31067431464183e+17, 1.31067431468558e+17, 1.310674314726205e+17, 1.310674314769955e+17, 1.31067431481058e+17, 1.31067431485433e+17, 1.310674314896518e+17, 1.310674314938705e+17, 1.310674314979329e+17, 1.310674315019955e+17, 1.310674315059018e+17, 1.310674315099643e+17, 1.310674315143392e+17, 1.310674315187142e+17, 1.310674315230893e+17, 1.310674315271517e+17, 1.310674315312142e+17, 1.31067431535433e+17, 1.310674315393393e+17, 1.310674315434017e+17, 1.310674315474642e+17, 1.310674315515268e+17, 1.310674315555892e+17, 1.310674315596517e+17, 1.310674315638705e+17, 1.310674315685581e+17, 1.310674315730893e+17, 1.310674315771517e+17, 1.310674315812142e+17, 1.31067431585433e+17, 1.310674315894956e+17, 1.310674315937142e+17, 1.310674315977768e+17, 1.310674316019955e+17, 1.31067431606058e+17, 1.310674316101204e+17, 1.310674316146518e+17, 1.310674316187142e+17, 1.310674316227768e+17, 1.310674316269955e+17, 1.310674316309016e+17, 1.310674316349642e+17, 1.310674316390268e+17, 1.310674316430893e+17, 1.310674316476205e+17, 1.310674316516829e+17, 1.310674316560581e+17, 1.310674316601204e+17, 1.310674316648079e+17, 1.310674316693393e+17, 1.310674316732454e+17, 1.31067431677308e+17, 1.310674316816829e+17, 1.310674316857455e+17, 1.310674316899643e+17, 1.310674316943393e+17, 1.310674316984017e+17, 1.310674317024643e+17, 1.310674317065267e+17, 1.310674317105892e+17, 1.310674317146518e+17, 1.310674317187142e+17, 1.310674317227767e+17, 1.310674317269955e+17, 1.31067431731058e+17, 1.310674317351205e+17, 1.31067431739183e+17, 1.310674317432454e+17, 1.310674317474642e+17, 1.310674317519955e+17, 1.31067431756058e+17, 1.310674317599643e+17, 1.31067431764183e+17, 1.31067431768558e+17, 1.310674317727768e+17, 1.310674317768393e+17, 1.310674317807455e+17, 1.310674317851205e+17, 1.310674317891831e+17, 1.310674317932456e+17, 1.310674317974642e+17, 1.310674318019955e+17, 1.310674318063704e+17, 1.31067431810433e+17, 1.310674318144955e+17, 1.31067431819183e+17, 1.310674318232456e+17, 1.31067431827308e+17, 1.310674318316831e+17, 1.310674318355892e+17, 1.310674318396517e+17, 1.310674318440268e+17, 1.310674318485581e+17, 1.310674318527767e+17, 1.310674318568393e+17, 1.310674318612142e+17, 1.31067431866058e+17, 1.310674318701204e+17, 1.31067431874183e+17, 1.310674318784018e+17, 1.310674318824643e+17, 1.310674318865267e+17, 1.31067431890433e+17, 1.310674318944955e+17, 1.310674318985581e+17, 1.310674319026205e+17, 1.31067431906683e+17, 1.310674319107455e+17, 1.310674319148081e+17, 1.310674319190268e+17, 1.310674319230892e+17, 1.310674319271517e+17, 1.310674319316829e+17, 1.310674319357455e+17, 1.310674319399643e+17, 1.310674319440268e+17, 1.310674319482455e+17, 1.31067431952308e+17, 1.310674319568393e+17, 1.310674319609018e+17, 1.31067431965433e+17, 1.310674319701206e+17, 1.31067431974183e+17, 1.310674319782455e+17, 1.31067431982308e+17, 1.310674319863704e+17, 1.31067431990433e+17, 1.310674319944955e+17, 1.31067431998558e+17, 1.310674320027767e+17, 1.310674320068393e+17, 1.310674320109018e+17, 1.310674320151205e+17, 1.31067432019183e+17, 1.310674320232456e+17, 1.31067432027308e+17, 1.310674320315268e+17, 1.310674320355892e+17, 1.310674320394956e+17, 1.31067432043558e+17, 1.310674320479331e+17, 1.310674320519955e+17, 1.31067432056058e+17, 1.310674320601204e+17, 1.31067432064183e+17, 1.310674320682455e+17, 1.310674320727768e+17, 1.310674320768392e+17, 1.310674320809018e+17, 1.310674320849642e+17, 1.310674320890267e+17, 1.310674320940268e+17, 1.310674320982455e+17, 1.310674321026205e+17, 1.310674321068393e+17, 1.310674321109018e+17, 1.310674321152768e+17, 1.310674321193393e+17, 1.310674321234017e+17, 1.310674321280893e+17, 1.310674321321517e+17, 1.31067432136058e+17, 1.31067432140433e+17, 1.310674321444956e+17, 1.310674321487142e+17, 1.31067432153558e+17, 1.310674321579331e+17, 1.310674321621518e+17, 1.310674321662143e+17, 1.310674321702767e+17, 1.310674321744955e+17, 1.310674321785581e+17, 1.310674321830892e+17, 1.310674321876205e+17, 1.310674321921517e+17, 1.310674321962143e+17, 1.310674322005892e+17, 1.310674322046518e+17, 1.310674322088705e+17, 1.31067432212933e+17, 1.310674322176205e+17, 1.310674322216831e+17, 1.31067432226058e+17, 1.31067432230433e+17, 1.310674322346518e+17, 1.310674322387142e+17, 1.310674322430893e+17, 1.310674322474642e+17, 1.310674322519955e+17, 1.31067432256058e+17, 1.310674322599643e+17, 1.310674322643392e+17, 1.310674322684018e+17, 1.310674322724643e+17, 1.310674322765267e+17, 1.310674322805893e+17, 1.310674322846516e+17, 1.31067432289183e+17, 1.310674322938706e+17, 1.310674322980892e+17, 1.310674323021517e+17, 1.310674323062143e+17, 1.310674323102767e+17, 1.310674323143392e+17, 1.31067432319183e+17, 1.310674323237143e+17, 1.310674323277768e+17, 1.310674323319954e+17, 1.31067432336058e+17, 1.310674323402767e+17, 1.310674323449642e+17, 1.310674323490267e+17, 1.310674323530893e+17, 1.310674323571517e+17, 1.310674323612142e+17, 1.31067432369183e+17, 1.310674323734017e+17, 1.310674323774642e+17, 1.310674323815268e+17, 1.31067432386058e+17, 1.310674323901204e+17, 1.31067432394183e+17, 1.31067432398558e+17, 1.310674324026205e+17, 1.31067432406683e+17, 1.31067432411058e+17, 1.310674324151205e+17, 1.310674324191831e+17, 1.310674324232456e+17, 1.310674324273079e+17, 1.310674324313705e+17, 1.310674324354331e+17, 1.310674324393393e+17, 1.310674324440268e+17, 1.310674324484018e+17, 1.310674324526205e+17, 1.31067432457308e+17, 1.310674324613705e+17, 1.310674324654331e+17, 1.310674324694956e+17, 1.310674324737143e+17, 1.310674324782455e+17, 1.310674324823081e+17, 1.310674324863704e+17, 1.310674324910579e+17, 1.310674324951205e+17, 1.310674324993393e+17, 1.310674325037143e+17, 1.310674325077768e+17, 1.310674325118392e+17, 1.310674325159017e+17, 1.310674325199643e+17, 1.310674325240268e+17, 1.310674325280892e+17, 1.310674325321517e+17, 1.310674325363706e+17, 1.310674325407455e+17, 1.310674325449642e+17, 1.31067432549183e+17, 1.310674325532456e+17, 1.31067432557308e+17, 1.310674325612143e+17, 1.310674325652767e+17, 1.310674325701204e+17, 1.310674325743392e+17, 1.31067432578558e+17, 1.310674325826205e+17, 1.310674325865267e+17, 1.31067432591058e+17, 1.310674325952768e+17, 1.310674325994956e+17, 1.310674326040268e+17, 1.310674326080893e+17, 1.310674326121518e+17, 1.310674326162143e+17, 1.310674326202767e+17, 1.310674326243393e+17, 1.310674326284017e+17, 1.310674326327767e+17, 1.310674326368393e+17, 1.310674326409018e+17, 1.310674326449642e+17, 1.310674326493393e+17, 1.310674326534017e+17, 1.310674326574642e+17, 1.310674326615268e+17, 1.310674326655892e+17, 1.310674326696517e+17, 1.310674326743392e+17, 1.310674326784018e+17, 1.310674326824643e+17, 1.310674326865267e+17, 1.31067432690433e+17, 1.310674326946516e+17, 1.31067432699183e+17, 1.31067432703558e+17, 1.310674327076205e+17, 1.310674327116829e+17, 1.310674327163704e+17, 1.31067432720433e+17, 1.310674327248081e+17, 1.310674327293393e+17, 1.310674327334017e+17, 1.310674327374643e+17, 1.310674327416831e+17, 1.310674327463704e+17, 1.310674327509018e+17, 1.31067432755433e+17, 1.310674327594954e+17, 1.31067432763558e+17, 1.310674327677768e+17, 1.310674327718392e+17, 1.310674327759017e+17, 1.310674327799643e+17, 1.310674327840268e+17, 1.310674327879331e+17, 1.310674327919955e+17, 1.310674327977768e+17, 1.310674328019955e+17, 1.310674328060581e+17, 1.310674328101204e+17, 1.310674328144955e+17, 1.31067432818558e+17, 1.31067432822933e+17, 1.31067432827308e+17, 1.310674328313705e+17, 1.31067432835433e+17, 1.310674328399643e+17, 1.310674328440268e+17, 1.310674328480892e+17, 1.310674328521518e+17, 1.310674328565267e+17, 1.31067432860433e+17, 1.310674328648079e+17, 1.310674328688704e+17, 1.31067432872933e+17, 1.31067432877308e+17, 1.310674328813705e+17, 1.31067432885433e+17, 1.310674328894956e+17, 1.31067432893558e+17, 1.310674328977768e+17, 1.310674329019955e+17, 1.310674329065267e+17, 1.310674329113705e+17, 1.310674329154331e+17, 1.310674329194954e+17, 1.31067432923558e+17, 1.310674329274643e+17, 1.310674329321517e+17, 1.310674329362143e+17, 1.31067432940433e+17, 1.310674329444955e+17, 1.310674329488705e+17, 1.31067432952933e+17, 1.310674329571517e+17, 1.310674329612142e+17, 1.310674329657455e+17, 1.31067432969808e+17, 1.310674329738705e+17, 1.310674329779331e+17, 1.310674329819955e+17, 1.31067432986058e+17, 1.310674329901204e+17, 1.310674329941829e+17, 1.310674329982455e+17, 1.310674330023081e+17, 1.310674330065267e+17},
			             {1.310674330065267e+17, 1.310674330109018e+17, 1.310674330149642e+17, 1.310674330190267e+17, 1.31067433023558e+17, 1.310674330276205e+17, 1.310674330316831e+17, 1.310674330359017e+17, 1.310674330399643e+17, 1.310674330438705e+17, 1.310674330482455e+17, 1.31067433052308e+17, 1.31067433056683e+17, 1.310674330609018e+17, 1.310674330654331e+17, 1.310674330699643e+17, 1.310674330740268e+17, 1.310674330780892e+17, 1.310674330824643e+17, 1.310674330865267e+17, 1.310674330905892e+17, 1.310674330946518e+17, 1.310674330987142e+17, 1.310674331027767e+17, 1.310674331068393e+17, 1.310674331107455e+17, 1.310674331151205e+17, 1.310674331193391e+17, 1.310674331232456e+17, 1.31067433127308e+17, 1.310674331316831e+17, 1.310674331357454e+17, 1.310674331399643e+17, 1.310674331443392e+17, 1.310674331484017e+17, 1.310674331524643e+17, 1.31067433156683e+17, 1.310674331607455e+17, 1.310674331649642e+17, 1.310674331694956e+17, 1.31067433173558e+17, 1.310674331777768e+17, 1.310674331821518e+17, 1.310674331862143e+17, 1.310674331902767e+17, 1.310674331948081e+17, 1.310674331988704e+17, 1.310674332034017e+17, 1.310674332074642e+17, 1.310674332121517e+17, 1.310674332165267e+17, 1.310674332207455e+17, 1.310674332249642e+17, 1.31067433229183e+17, 1.310674332334017e+17, 1.310674332374643e+17, 1.310674332416831e+17, 1.310674332459018e+17, 1.310674332499642e+17, 1.310674332541829e+17, 1.310674332582455e+17, 1.310674332624643e+17, 1.310674332665268e+17, 1.310674332705892e+17, 1.310674332746518e+17, 1.31067433278558e+17, 1.31067433282933e+17, 1.310674332869955e+17, 1.310674332909018e+17, 1.310674332951205e+17, 1.31067433299183e+17, 1.310674333030893e+17, 1.310674333076205e+17, 1.310674333118392e+17, 1.310674333159017e+17, 1.310674333201204e+17, 1.310674333243393e+17, 1.310674333288705e+17, 1.31067433332933e+17, 1.310674333369956e+17, 1.310674333409018e+17, 1.310674333449642e+17, 1.310674333490267e+17, 1.310674333532454e+17, 1.31067433357308e+17, 1.310674333613705e+17, 1.310674333657455e+17, 1.31067433369808e+17, 1.310674333738705e+17, 1.310674333780892e+17, 1.310674333824643e+17, 1.310674333868393e+17, 1.310674333909018e+17, 1.310674333951204e+17, 1.310674333993393e+17, 1.310674334034017e+17, 1.310674334076205e+17, 1.310674334116831e+17, 1.310674334159018e+17, 1.31067433420433e+17, 1.310674334244955e+17, 1.31067433428558e+17, 1.310674334326205e+17, 1.31067433436683e+17, 1.310674334409018e+17, 1.31067433445433e+17, 1.310674334494956e+17, 1.31067433453558e+17, 1.310674334579331e+17, 1.310674334619955e+17, 1.31067433466058e+17, 1.310674334701204e+17, 1.31067433474183e+17, 1.310674334784017e+17, 1.310674334824643e+17, 1.310674334865267e+17, 1.310674334909018e+17, 1.310674334949642e+17, 1.310674334990267e+17, 1.310674335038705e+17, 1.310674335082455e+17, 1.310674335130893e+17, 1.310674335171517e+17, 1.310674335212143e+17, 1.310674335252768e+17, 1.310674335293393e+17, 1.310674335334017e+17, 1.310674335374643e+17, 1.310674335415268e+17, 1.310674335455892e+17, 1.310674335499643e+17, 1.310674335540268e+17, 1.310674335580893e+17, 1.310674335619955e+17, 1.310674335662143e+17, 1.310674335701204e+17, 1.31067433574183e+17, 1.310674335782455e+17, 1.310674335824643e+17, 1.31067433586683e+17, 1.310674335907455e+17, 1.310674335949642e+17, 1.310674335990268e+17, 1.310674336030893e+17, 1.310674336071516e+17, 1.310674336118392e+17, 1.310674336159018e+17, 1.310674336199642e+17, 1.310674336240268e+17, 1.310674336280892e+17, 1.310674336321518e+17, 1.310674336371517e+17, 1.310674336413705e+17, 1.310674336455892e+17, 1.310674336502767e+17, 1.310674336543393e+17, 1.310674336582455e+17, 1.31067433662308e+17, 1.31067433666683e+17, 1.310674336707455e+17, 1.310674336748081e+17, 1.310674336787142e+17, 1.310674336830893e+17, 1.310674336874643e+17, 1.310674336915268e+17, 1.310674336960581e+17, 1.310674337002767e+17, 1.310674337043392e+17, 1.310674337090268e+17, 1.310674337132454e+17, 1.31067433717308e+17, 1.310674337212142e+17, 1.310674337255892e+17, 1.31067433729808e+17, 1.310674337338705e+17, 1.310674337380892e+17, 1.310674337423081e+17, 1.310674337463706e+17, 1.31067433750433e+17, 1.310674337549642e+17, 1.310674337590267e+17, 1.310674337630893e+17, 1.310674337671517e+17, 1.310674337712142e+17, 1.310674337752767e+17, 1.310674337794956e+17, 1.310674337840268e+17, 1.310674337882455e+17, 1.31067433792308e+17, 1.310674337963706e+17, 1.310674338005893e+17, 1.310674338046518e+17, 1.310674338090268e+17, 1.310674338132456e+17, 1.31067433817308e+17, 1.310674338213705e+17, 1.310674338254331e+17, 1.310674338294954e+17, 1.31067433833558e+17, 1.310674338376205e+17, 1.310674338419955e+17, 1.310674338460581e+17, 1.310674338505893e+17, 1.310674338546518e+17, 1.310674338590268e+17, 1.31067433863558e+17, 1.310674338685581e+17, 1.310674338726204e+17, 1.310674338768392e+17, 1.310674338809018e+17, 1.310674338848079e+17, 1.310674338890267e+17, 1.310674338930893e+17, 1.310674338971517e+17, 1.310674339015268e+17, 1.310674339057455e+17, 1.31067433909808e+17, 1.310674339138705e+17, 1.310674339180892e+17, 1.310674339221518e+17, 1.310674339262143e+17, 1.310674339302767e+17, 1.310674339343392e+17, 1.310674339384018e+17, 1.310674339424643e+17, 1.310674339465267e+17, 1.310674339516829e+17, 1.310674339557454e+17, 1.31067433959808e+17, 1.310674339640268e+17, 1.310674339679331e+17, 1.310674339719955e+17, 1.310674339765267e+17, 1.310674339807455e+17, 1.310674339848081e+17, 1.310674339888705e+17, 1.310674339932456e+17, 1.31067433997308e+17, 1.310674340013705e+17, 1.31067434005433e+17, 1.310674340094956e+17, 1.310674340134017e+17, 1.310674340176205e+17, 1.310674340215268e+17, 1.310674340257454e+17, 1.31067434029808e+17, 1.310674340338706e+17, 1.310674340379329e+17, 1.310674340419955e+17, 1.31067434046058e+17, 1.310674340501204e+17, 1.31067434054183e+17, 1.310674340582455e+17, 1.310674340623081e+17, 1.310674340663704e+17, 1.310674340709018e+17, 1.310674340749642e+17, 1.310674340790268e+17, 1.310674340830893e+17, 1.31067434087308e+17, 1.310674340913705e+17, 1.310674340952768e+17, 1.310674340993393e+17, 1.310674341037143e+17, 1.310674341077768e+17, 1.310674341121518e+17, 1.310674341168392e+17, 1.310674341210579e+17, 1.31067434125433e+17, 1.310674341294954e+17, 1.31067434133558e+17, 1.310674341379329e+17, 1.310674341419955e+17, 1.31067434146058e+17, 1.310674341505893e+17, 1.310674341546518e+17, 1.310674341587142e+17, 1.310674341627767e+17, 1.310674341668393e+17, 1.310674341707455e+17, 1.310674341748081e+17, 1.310674341790268e+17, 1.310674341830892e+17, 1.310674341871517e+17, 1.31067434191058e+17, 1.31067434196058e+17, 1.310674342001204e+17, 1.31067434204183e+17, 1.310674342082455e+17, 1.310674342124643e+17, 1.310674342168393e+17, 1.31067434221058e+17, 1.31067434225433e+17, 1.31067434229808e+17, 1.310674342340268e+17, 1.310674342380893e+17, 1.310674342426204e+17, 1.310674342468392e+17, 1.310674342515268e+17, 1.310674342555892e+17, 1.31067434259808e+17, 1.310674342638705e+17, 1.310674342680892e+17, 1.310674342724643e+17, 1.310674342765267e+17, 1.310674342805893e+17, 1.310674342846518e+17, 1.310674342887142e+17, 1.310674342927768e+17, 1.310674342969955e+17, 1.31067434301058e+17, 1.310674343051205e+17, 1.310674343096518e+17, 1.310674343137142e+17, 1.310674343177768e+17, 1.310674343219955e+17, 1.310674343260581e+17, 1.310674343301204e+17, 1.31067434334183e+17, 1.310674343384018e+17, 1.310674343424643e+17, 1.31067434346683e+17, 1.310674343507455e+17, 1.310674343549642e+17, 1.310674343590267e+17, 1.310674343630893e+17, 1.310674343671517e+17, 1.310674343712142e+17, 1.310674343752768e+17, 1.310674343793393e+17, 1.310674343834017e+17, 1.310674343876205e+17, 1.310674343916831e+17, 1.310674343957454e+17, 1.310674344002767e+17, 1.310674344043393e+17, 1.31067434408558e+17, 1.310674344126204e+17, 1.310674344165268e+17, 1.310674344205892e+17, 1.310674344248079e+17, 1.310674344288705e+17, 1.31067434433558e+17, 1.310674344374642e+17, 1.310674344419955e+17, 1.31067434446058e+17, 1.310674344502767e+17, 1.310674344546516e+17, 1.310674344587142e+17, 1.310674344630893e+17, 1.310674344671517e+17, 1.310674344712143e+17, 1.310674344754331e+17, 1.31067434479808e+17, 1.310674344838705e+17, 1.310674344879331e+17, 1.310674344924643e+17, 1.310674344965267e+17, 1.310674345005892e+17, 1.310674345054331e+17, 1.310674345094956e+17, 1.310674345141829e+17, 1.310674345182455e+17, 1.310674345223081e+17, 1.310674345265267e+17, 1.310674345305892e+17, 1.310674345346518e+17, 1.310674345387142e+17, 1.310674345432454e+17, 1.31067434547308e+17, 1.310674345513705e+17, 1.310674345559017e+17, 1.310674345599643e+17, 1.310674345640268e+17, 1.310674345680892e+17, 1.310674345721517e+17, 1.310674345762143e+17, 1.31067434580433e+17, 1.310674345848081e+17, 1.310674345888704e+17, 1.310674345934017e+17, 1.310674345980892e+17, 1.310674346019955e+17, 1.310674346068393e+17, 1.310674346112142e+17, 1.31067434615433e+17, 1.310674346194956e+17, 1.31067434623558e+17, 1.310674346280892e+17, 1.310674346321518e+17, 1.310674346363706e+17, 1.310674346443393e+17, 1.310674346490267e+17, 1.310674346530893e+17, 1.310674346571517e+17, 1.310674346613705e+17, 1.31067434665433e+17, 1.310674346694956e+17, 1.310674346743392e+17, 1.310674346787142e+17, 1.310674346827767e+17, 1.310674346873079e+17, 1.310674346915268e+17, 1.310674346957454e+17, 1.310674346999643e+17, 1.310674347040268e+17, 1.310674347080893e+17, 1.310674347124643e+17, 1.310674347163704e+17, 1.31067434720433e+17, 1.310674347244955e+17, 1.31067434728558e+17, 1.310674347326205e+17, 1.31067434736683e+17, 1.310674347407455e+17, 1.310674347448079e+17, 1.310674347488705e+17, 1.31067434753558e+17, 1.310674347576205e+17, 1.310674347618392e+17, 1.310674347659018e+17, 1.310674347702767e+17, 1.310674347743393e+17, 1.310674347787142e+17, 1.310674347830893e+17, 1.31067434787308e+17, 1.310674347913705e+17, 1.31067434795433e+17, 1.310674347994954e+17, 1.31067434803558e+17, 1.310674348076205e+17, 1.310674348116831e+17, 1.310674348157455e+17, 1.310674348202767e+17, 1.310674348243392e+17, 1.310674348284018e+17, 1.310674348330893e+17, 1.310674348373079e+17, 1.310674348413705e+17, 1.310674348454331e+17, 1.310674348493393e+17, 1.310674348537142e+17, 1.310674348579331e+17, 1.310674348619955e+17, 1.31067434866058e+17, 1.310674348701204e+17, 1.310674348744955e+17, 1.310674348787142e+17, 1.310674348830893e+17, 1.310674348874643e+17, 1.310674348915268e+17, 1.310674348957455e+17, 1.310674349002767e+17, 1.310674349043393e+17, 1.310674349084017e+17, 1.310674349127767e+17, 1.310674349168392e+17, 1.310674349209018e+17, 1.31067434925433e+17, 1.310674349294956e+17, 1.31067434933558e+17, 1.310674349376205e+17, 1.310674349415268e+17, 1.310674349455892e+17, 1.310674349496517e+17, 1.310674349538705e+17, 1.310674349582455e+17, 1.31067434962308e+17, 1.310674349665267e+17, 1.310674349709016e+17, 1.310674349748081e+17, 1.310674349791831e+17, 1.310674349832454e+17, 1.310674349871517e+17, 1.310674349926205e+17, 1.31067434996683e+17, 1.310674350007455e+17, 1.310674350048079e+17, 1.310674350088705e+17, 1.310674350132456e+17, 1.310674350177766e+17, 1.310674350218392e+17, 1.310674350259018e+17, 1.310674350299642e+17, 1.310674350338705e+17, 1.310674350382455e+17, 1.310674350423081e+17, 1.310674350462143e+17, 1.310674350505892e+17, 1.310674350546518e+17, 1.310674350587144e+17, 1.310674350627767e+17, 1.31067435066683e+17, 1.310674350712142e+17, 1.31067435076058e+17, 1.310674350802767e+17, 1.310674350843392e+17, 1.310674350885581e+17, 1.310674350930893e+17, 1.310674350971517e+17, 1.310674351012143e+17, 1.310674351052767e+17, 1.310674351093393e+17, 1.31067435113558e+17, 1.310674351182455e+17, 1.31067435122308e+17, 1.310674351265267e+17, 1.310674351305892e+17, 1.310674351346518e+17, 1.310674351387142e+17, 1.31067435142933e+17, 1.310674351469955e+17, 1.31067435151058e+17, 1.31067435155433e+17, 1.310674351594956e+17, 1.310674351640268e+17, 1.310674351680893e+17, 1.31067435172308e+17, 1.310674351765268e+17, 1.310674351805892e+17, 1.310674351846518e+17, 1.310674351888705e+17, 1.310674351929331e+17, 1.310674351969955e+17, 1.31067435201058e+17, 1.31067435205433e+17, 1.310674352094956e+17, 1.31067435213558e+17, 1.310674352174642e+17, 1.310674352219955e+17, 1.31067435226058e+17, 1.310674352301206e+17, 1.310674352340268e+17, 1.310674352380892e+17, 1.310674352421518e+17, 1.310674352463706e+17, 1.310674352502767e+17, 1.310674352543393e+17, 1.310674352584017e+17, 1.310674352624643e+17, 1.31067435266683e+17, 1.310674352709018e+17, 1.310674352749642e+17, 1.310674352796517e+17, 1.310674352840268e+17, 1.310674352880892e+17, 1.310674352919955e+17, 1.31067435296058e+17, 1.310674353005893e+17, 1.310674353048081e+17, 1.310674353090268e+17, 1.310674353130893e+17, 1.310674353174643e+17, 1.310674353218392e+17, 1.310674353263704e+17, 1.31067435330433e+17, 1.310674353344956e+17, 1.310674353390268e+17, 1.310674353430893e+17, 1.310674353471517e+17, 1.310674353512142e+17, 1.310674353552768e+17, 1.310674353593393e+17, 1.310674353634017e+17, 1.310674353674642e+17, 1.310674353715268e+17, 1.31067435376058e+17, 1.310674353805893e+17, 1.310674353848081e+17, 1.310674353891831e+17, 1.310674353934017e+17, 1.310674353974642e+17, 1.310674354015268e+17, 1.310674354057455e+17, 1.310674354099643e+17, 1.31067435414183e+17, 1.310674354182455e+17, 1.31067435422308e+17, 1.310674354265267e+17, 1.310674354309018e+17, 1.310674354349642e+17, 1.310674354396517e+17, 1.310674354437142e+17, 1.310674354476205e+17, 1.310674354516831e+17, 1.310674354565267e+17, 1.310674354609018e+17, 1.31067435465433e+17, 1.310674354693393e+17, 1.310674354740268e+17, 1.310674354780892e+17, 1.310674354824643e+17, 1.31067435487308e+17, 1.310674354916829e+17, 1.310674354959017e+17, 1.310674355001204e+17, 1.31067435504183e+17, 1.310674355080892e+17, 1.310674355121517e+17, 1.310674355162143e+17, 1.310674355202767e+17, 1.310674355243392e+17, 1.310674355284018e+17, 1.310674355324643e+17, 1.310674355363706e+17, 1.310674355407455e+17, 1.310674355451204e+17, 1.31067435549183e+17, 1.310674355534017e+17, 1.310674355574643e+17, 1.310674355615267e+17, 1.31067435565433e+17, 1.310674355694956e+17, 1.310674355737142e+17, 1.310674355777768e+17, 1.310674355818392e+17, 1.310674355859017e+17, 1.310674355899643e+17, 1.310674355940268e+17, 1.310674355982455e+17, 1.31067435602308e+17, 1.310674356062143e+17, 1.310674356112142e+17, 1.31067435615433e+17, 1.31067435619808e+17, 1.310674356240268e+17, 1.310674356282455e+17, 1.310674356323081e+17, 1.310674356363706e+17, 1.310674356404329e+17, 1.310674356444955e+17, 1.310674356485581e+17, 1.310674356526204e+17, 1.31067435656683e+17, 1.310674356607455e+17, 1.310674356652767e+17, 1.310674356693393e+17, 1.310674356734017e+17, 1.310674356774642e+17, 1.310674356815268e+17, 1.31067435685433e+17, 1.310674356894954e+17, 1.310674356940268e+17, 1.31067435698558e+17, 1.31067435702933e+17, 1.31067435707308e+17, 1.310674357113705e+17, 1.310674357155892e+17, 1.310674357196518e+17, 1.310674357237142e+17, 1.310674357276205e+17, 1.310674357321517e+17, 1.310674357362143e+17, 1.310674357402767e+17, 1.310674357444955e+17, 1.31067435748558e+17, 1.310674357532454e+17, 1.31067435757308e+17, 1.310674357618392e+17, 1.310674357662141e+17, 1.310674357702767e+17, 1.310674357743393e+17, 1.310674357784017e+17, 1.310674357824643e+17, 1.310674357868393e+17, 1.310674357913705e+17, 1.31067435796058e+17, 1.310674358009018e+17, 1.310674358049642e+17, 1.310674358090268e+17, 1.310674358130893e+17, 1.310674358171517e+17, 1.310674358212143e+17, 1.310674358252768e+17, 1.310674358293393e+17, 1.310674358334017e+17, 1.310674358374643e+17, 1.310674358415268e+17, 1.310674358459017e+17, 1.310674358499643e+17, 1.310674358540268e+17, 1.310674358579329e+17, 1.310674358621517e+17, 1.31067435866058e+17, 1.310674358701204e+17, 1.31067435874183e+17, 1.310674358782455e+17, 1.31067435882308e+17, 1.310674358863704e+17, 1.31067435890433e+17, 1.310674358944955e+17, 1.31067435898558e+17, 1.310674359026205e+17, 1.31067435906683e+17, 1.310674359107455e+17, 1.310674359148081e+17, 1.310674359188705e+17, 1.310674359230893e+17, 1.310674359271517e+17, 1.310674359312143e+17, 1.310674359352768e+17, 1.310674359393393e+17, 1.310674359432456e+17, 1.310674359480893e+17, 1.310674359521517e+17, 1.31067435956058e+17, 1.310674359601204e+17, 1.310674359641829e+17, 1.310674359682455e+17, 1.310674359723081e+17, 1.310674359763704e+17, 1.310674359807455e+17, 1.310674359848081e+17, 1.310674359888705e+17, 1.310674359930893e+17, 1.310674359971517e+17, 1.310674360012142e+17, 1.310674360051205e+17, 1.310674360094956e+17, 1.31067436013558e+17, 1.310674360176205e+17, 1.310674360216831e+17, 1.31067436026058e+17, 1.310674360301204e+17, 1.310674360341829e+17, 1.310674360387142e+17, 1.310674360427768e+17, 1.310674360468393e+17, 1.310674360513705e+17, 1.31067436055433e+17, 1.310674360596517e+17, 1.310674360637143e+17, 1.310674360679331e+17, 1.31067436072933e+17, 1.310674360769955e+17, 1.31067436081058e+17, 1.310674360852768e+17, 1.310674360893393e+17, 1.310674360937142e+17, 1.310674360977768e+17, 1.310674361018392e+17, 1.310674361057454e+17, 1.31067436109808e+17, 1.310674361138706e+17, 1.310674361180892e+17, 1.310674361221517e+17, 1.310674361262143e+17, 1.310674361307455e+17, 1.310674361349642e+17, 1.310674361390267e+17, 1.31067436142933e+17, 1.310674361469955e+17, 1.31067436151058e+17, 1.310674361551205e+17, 1.310674361596517e+17, 1.310674361637143e+17, 1.310674361677766e+17, 1.310674361718392e+17, 1.310674361759018e+17, 1.310674361799643e+17, 1.310674361840268e+17, 1.310674361884017e+17, 1.310674361924643e+17, 1.310674361965268e+17, 1.310674362005892e+17, 1.310674362046518e+17, 1.310674362087144e+17, 1.310674362127767e+17, 1.310674362168392e+17, 1.310674362212142e+17, 1.310674362252768e+17, 1.310674362293393e+17, 1.31067436233558e+17, 1.310674362379331e+17, 1.310674362419955e+17, 1.31067436246058e+17, 1.31067436250433e+17, 1.310674362546516e+17, 1.310674362588705e+17, 1.31067436262933e+17, 1.310674362674642e+17, 1.310674362715268e+17, 1.310674362755892e+17, 1.310674362799643e+17, 1.31067436284183e+17, 1.310674362880892e+17, 1.310674362924643e+17, 1.310674362969955e+17, 1.31067436301058e+17, 1.310674363055892e+17, 1.31067436309808e+17, 1.310674363143393e+17, 1.310674363184017e+17, 1.310674363224643e+17, 1.310674363265268e+17, 1.310674363309018e+17, 1.310674363349642e+17, 1.31067436339183e+17, 1.310674363432454e+17, 1.31067436347308e+17, 1.310674363513705e+17, 1.31067436355433e+17, 1.310674363601204e+17, 1.31067436364183e+17, 1.310674363680892e+17, 1.310674363721518e+17, 1.310674363765267e+17, 1.310674363805893e+17, 1.310674363846516e+17, 1.310674363887142e+17, 1.310674363927768e+17, 1.310674363968392e+17, 1.310674364007455e+17, 1.310674364048079e+17, 1.310674364099643e+17, 1.31067436414183e+17, 1.310674364187142e+17, 1.310674364227767e+17, 1.310674364269956e+17, 1.310674364315268e+17, 1.310674364355892e+17, 1.310674364396517e+17, 1.310674364437143e+17, 1.310674364476205e+17, 1.310674364518392e+17, 1.310674364559018e+17, 1.310674364602767e+17, 1.310674364643392e+17, 1.310674364687144e+17, 1.310674364727767e+17, 1.310674364771517e+17, 1.310674364813705e+17, 1.310674364857455e+17, 1.31067436489808e+17, 1.310674364938705e+17, 1.310674364980892e+17, 1.310674365024643e+17, 1.310674365065267e+17, 1.310674365109018e+17, 1.310674365149644e+17, 1.310674365190268e+17, 1.310674365230893e+17, 1.310674365271517e+17, 1.310674365312143e+17, 1.310674365362143e+17, 1.31067436540433e+17, 1.310674365446518e+17, 1.310674365488705e+17, 1.310674365532456e+17, 1.310674365574643e+17, 1.310674365616831e+17, 1.310674365659018e+17, 1.310674365699642e+17, 1.310674365740268e+17, 1.310674365782455e+17, 1.310674365823081e+17, 1.31067436586683e+17, 1.310674365909018e+17, 1.310674365949642e+17, 1.310674365990267e+17, 1.310674366032454e+17, 1.31067436607308e+17, 1.310674366116829e+17, 1.310674366159017e+17, 1.310674366199643e+17, 1.310674366243393e+17, 1.310674366284018e+17, 1.310674366327768e+17, 1.31067436637308e+17, 1.310674366413705e+17, 1.310674366459017e+17, 1.310674366502767e+17, 1.310674366543392e+17, 1.310674366588705e+17, 1.310674366632456e+17, 1.310674366674643e+17, 1.310674366716831e+17, 1.310674366757455e+17, 1.31067436679808e+17, 1.310674366838705e+17, 1.310674366879331e+17, 1.310674366919955e+17, 1.31067436696058e+17, 1.310674367001206e+17, 1.310674367044955e+17, 1.31067436708558e+17, 1.310674367126204e+17, 1.310674367169955e+17, 1.310674367210579e+17, 1.310674367257455e+17, 1.310674367299643e+17, 1.310674367340268e+17, 1.310674367382455e+17, 1.310674367427768e+17, 1.310674367468393e+17, 1.310674367512143e+17, 1.310674367555892e+17, 1.310674367596518e+17, 1.310674367638705e+17, 1.310674367679329e+17, 1.310674367724643e+17, 1.310674367768393e+17, 1.310674367809018e+17, 1.310674367849642e+17, 1.310674367890268e+17, 1.310674367930893e+17, 1.310674367977766e+17, 1.310674368018392e+17, 1.31067436806058e+17, 1.310674368101204e+17, 1.310674368141829e+17, 1.310674368188705e+17, 1.31067436822933e+17, 1.310674368269955e+17, 1.310674368313705e+17, 1.31067436835433e+17, 1.310674368394956e+17, 1.310674368434017e+17, 1.310674368474642e+17, 1.310674368516831e+17, 1.310674368559017e+17, 1.310674368601204e+17, 1.310674368644955e+17, 1.310674368687142e+17, 1.310674368727767e+17, 1.310674368771517e+17, 1.310674368812143e+17, 1.310674368852767e+17, 1.310674368893393e+17, 1.310674368937142e+17, 1.310674368979331e+17, 1.310674369019955e+17, 1.31067436906058e+17, 1.310674369101204e+17, 1.31067436914183e+17, 1.310674369182456e+17, 1.310674369224643e+17, 1.310674369265267e+17, 1.310674369305893e+17, 1.310674369346518e+17, 1.310674369387142e+17, 1.31067436942933e+17, 1.310674369469956e+17, 1.31067436951058e+17, 1.310674369559018e+17, 1.31067436959808e+17, 1.310674369640268e+17, 1.310674369680893e+17, 1.310674369721517e+17, 1.310674369762143e+17, 1.310674369807455e+17, 1.310674369849642e+17, 1.310674369896517e+17, 1.310674369937143e+17, 1.310674369979331e+17, 1.310674370021518e+17, 1.310674370062143e+17, 1.310674370104329e+17, 1.310674370144955e+17, 1.310674370184018e+17, 1.310674370265268e+17, 1.310674370305893e+17, 1.310674370344955e+17, 1.310674370387142e+17, 1.310674370427768e+17, 1.310674370468392e+17, 1.310674370510579e+17, 1.31067437055433e+17, 1.310674370596517e+17, 1.310674370637143e+17, 1.310674370680892e+17, 1.310674370724643e+17, 1.310674370765267e+17, 1.310674370809018e+17, 1.310674370851205e+17, 1.310674370894956e+17, 1.310674370940268e+17, 1.310674370987144e+17, 1.31067437102933e+17, 1.310674371069955e+17, 1.31067437111058e+17, 1.310674371149642e+17, 1.310674371190268e+17, 1.310674371230893e+17, 1.310674371271517e+17, 1.310674371312142e+17, 1.31067437136058e+17, 1.310674371401204e+17, 1.310674371440268e+17, 1.310674371484018e+17, 1.310674371524643e+17, 1.31067437156683e+17, 1.310674371613705e+17, 1.310674371659017e+17, 1.310674371702767e+17, 1.310674371743392e+17, 1.310674371784018e+17, 1.310674371824643e+17, 1.310674371865267e+17, 1.310674371905893e+17, 1.310674371944955e+17, 1.310674371988705e+17, 1.31067437202933e+17, 1.310674372074643e+17, 1.310674372115268e+17, 1.310674372154331e+17, 1.310674372194956e+17, 1.310674372237142e+17, 1.310674372280893e+17, 1.310674372321517e+17, 1.310674372362143e+17, 1.31067437240433e+17, 1.310674372444955e+17, 1.31067437248558e+17, 1.310674372526205e+17, 1.310674372569955e+17, 1.31067437261058e+17, 1.310674372649642e+17, 1.31067437269808e+17, 1.31067437274183e+17, 1.310674372782455e+17, 1.31067437282308e+17, 1.310674372863706e+17, 1.31067437290433e+17, 1.310674372944955e+17, 1.310674372985581e+17, 1.310674373024643e+17, 1.310674373065267e+17, 1.310674373105892e+17, 1.310674373151205e+17, 1.310674373193393e+17, 1.310674373234017e+17, 1.310674373274642e+17, 1.310674373316829e+17, 1.310674373357455e+17, 1.31067437339808e+17, 1.310674373440268e+17, 1.310674373480892e+17, 1.310674373521517e+17, 1.310674373562143e+17, 1.310674373602767e+17, 1.310674373643393e+17, 1.310674373684018e+17, 1.310674373724643e+17, 1.310674373768393e+17, 1.310674373809016e+17, 1.310674373848081e+17, 1.310674373899643e+17, 1.310674373943392e+17, 1.310674373990267e+17, 1.310674374030893e+17, 1.310674374071517e+17, 1.310674374113705e+17, 1.31067437415433e+17, 1.310674374193393e+17, 1.310674374238705e+17, 1.310674374279331e+17, 1.31067437432308e+17, 1.310674374363706e+17, 1.31067437440433e+17, 1.310674374444955e+17, 1.310674374484017e+17, 1.310674374526204e+17, 1.310674374568393e+17, 1.310674374609018e+17, 1.310674374649644e+17, 1.31067437469183e+17, 1.310674374732454e+17, 1.310674374771517e+17, 1.310674374812142e+17, 1.310674374857455e+17, 1.31067437489808e+17, 1.310674374938705e+17, 1.310674374977768e+17, 1.310674375019955e+17, 1.310674375063706e+17, 1.31067437510433e+17, 1.310674375144955e+17, 1.310674375185581e+17, 1.310674375227768e+17, 1.31067437527308e+17, 1.310674375315268e+17, 1.310674375359017e+17, 1.310674375401204e+17, 1.310674375443392e+17, 1.31067437548558e+17, 1.310674375526205e+17, 1.31067437556683e+17, 1.310674375609018e+17, 1.310674375652768e+17, 1.310674375693393e+17, 1.310674375734017e+17, 1.310674375774643e+17, 1.310674375821518e+17, 1.310674375862143e+17, 1.310674375901206e+17, 1.310674375982455e+17, 1.310674376023081e+17, 1.310674376062143e+17, 1.310674376102769e+17, 1.310674376149642e+17, 1.31067437619183e+17, 1.310674376232456e+17, 1.310674376276205e+17, 1.310674376321518e+17, 1.310674376365267e+17, 1.310674376405893e+17, 1.310674376448081e+17, 1.310674376490268e+17, 1.310674376530893e+17, 1.310674376573079e+17, 1.310674376616829e+17, 1.310674376657455e+17, 1.310674376701204e+17, 1.310674376749642e+17, 1.310674376790268e+17, 1.310674376834017e+17, 1.310674376874643e+17, 1.310674376918392e+17, 1.31067437696058e+17, 1.310674377002767e+17, 1.310674377043393e+17, 1.310674377084017e+17, 1.310674377124643e+17, 1.31067437716683e+17, 1.310674377210579e+17, 1.310674377255892e+17, 1.310674377301204e+17, 1.31067437734183e+17, 1.310674377382455e+17, 1.310674377426205e+17, 1.31067437746683e+17, 1.310674377507455e+17, 1.310674377546518e+17, 1.310674377587142e+17, 1.310674377627767e+17, 1.310674377668393e+17, 1.310674377707455e+17, 1.310674377748081e+17, 1.310674377788704e+17, 1.31067437782933e+17, 1.310674377869956e+17, 1.310674377910579e+17, 1.310674377951205e+17, 1.310674377996517e+17, 1.310674378037143e+17, 1.310674378077768e+17, 1.310674378119955e+17, 1.31067437816058e+17, 1.310674378201204e+17, 1.31067437824183e+17, 1.310674378280892e+17, 1.310674378321517e+17, 1.310674378362143e+17, 1.310674378402767e+17, 1.310674378443393e+17, 1.310674378482455e+17, 1.310674378526205e+17, 1.31067437856683e+17, 1.310674378607455e+17, 1.310674378649642e+17, 1.310674378693393e+17, 1.31067437873558e+17, 1.310674378776205e+17, 1.310674378815268e+17, 1.310674378859017e+17, 1.310674378899643e+17, 1.310674378940268e+17, 1.310674378980892e+17, 1.31067437902308e+17, 1.310674379063704e+17, 1.31067437910433e+17, 1.310674379148081e+17, 1.310674379188705e+17, 1.31067437922933e+17, 1.310674379271517e+17, 1.310674379312142e+17, 1.310674379352768e+17, 1.310674379393393e+17, 1.310674379434017e+17, 1.310674379474643e+17, 1.310674379515268e+17, 1.310674379554331e+17, 1.310674379596517e+17, 1.310674379637143e+17, 1.310674379677768e+17, 1.310674379718392e+17, 1.310674379759018e+17, 1.310674379799642e+17, 1.31067437984183e+17, 1.310674379880893e+17, 1.310674379921517e+17, 1.310674379962143e+17, 1.310674380002767e+17, 1.310674380043392e+17, 1.310674380084018e+17, 1.310674380124643e+17, 1.31067438017308e+17, 1.310674380213705e+17, 1.31067438025433e+17, 1.310674380296517e+17, 1.310674380338705e+17, 1.310674380377768e+17, 1.310674380419955e+17, 1.31067438046058e+17, 1.310674380501206e+17, 1.31067438054183e+17, 1.310674380582455e+17, 1.31067438063558e+17, 1.310674380676206e+17, 1.31067438072308e+17, 1.310674380763704e+17, 1.31067438080433e+17, 1.310674380844955e+17, 1.31067438088558e+17, 1.310674380926205e+17, 1.310674380971517e+17, 1.310674381015267e+17, 1.310674381059018e+17, 1.310674381102767e+17, 1.310674381144956e+17, 1.310674381190267e+17, 1.310674381230893e+17, 1.310674381269955e+17, 1.310674381312142e+17, 1.31067438135433e+17, 1.310674381394956e+17, 1.31067438144183e+17, 1.310674381482455e+17, 1.31067438152308e+17, 1.310674381563706e+17, 1.310674381602767e+17, 1.310674381643393e+17, 1.310674381688704e+17, 1.310674381730893e+17, 1.310674381779329e+17, 1.310674381824643e+17, 1.310674381865267e+17, 1.31067438191058e+17, 1.310674381951205e+17, 1.310674381993393e+17, 1.310674382034017e+17, 1.310674382076205e+17, 1.310674382116831e+17, 1.310674382159018e+17, 1.310674382201206e+17, 1.310674382246516e+17, 1.310674382288705e+17, 1.310674382334017e+17, 1.310674382376205e+17, 1.310674382416829e+17, 1.310674382457455e+17, 1.31067438249808e+17, 1.310674382538705e+17, 1.310674382582455e+17, 1.310674382626205e+17, 1.31067438266683e+17, 1.310674382705893e+17, 1.310674382748081e+17, 1.310674382790268e+17, 1.310674382832456e+17, 1.310674382877768e+17, 1.310674382919955e+17, 1.310674382960581e+17, 1.310674382999643e+17, 1.310674383046518e+17, 1.310674383087142e+17, 1.310674383127767e+17, 1.31067438317308e+17, 1.310674383218392e+17, 1.310674383262141e+17, 1.310674383302767e+17, 1.310674383343393e+17, 1.310674383385581e+17, 1.31067438342933e+17, 1.310674383479331e+17, 1.310674383519955e+17, 1.310674383562143e+17, 1.31067438360433e+17, 1.310674383644955e+17, 1.310674383687142e+17, 1.310674383730893e+17, 1.310674383774643e+17, 1.310674383819955e+17, 1.31067438386058e+17, 1.310674383901204e+17, 1.31067438394183e+17, 1.310674383982455e+17, 1.31067438402308e+17, 1.310674384063704e+17, 1.310674384102767e+17, 1.310674384143392e+17, 1.31067438418558e+17, 1.310674384226204e+17, 1.310674384269955e+17, 1.31067438431058e+17, 1.310674384349642e+17, 1.310674384390267e+17, 1.310674384430893e+17, 1.310674384471517e+17, 1.310674384512142e+17, 1.310674384552768e+17, 1.310674384593393e+17, 1.31067438463558e+17, 1.310674384676205e+17, 1.310674384719955e+17, 1.31067438476058e+17, 1.310674384805892e+17, 1.310674384851205e+17, 1.31067438489183e+17, 1.310674384932454e+17, 1.310674384971517e+17, 1.310674385013705e+17, 1.310674385057455e+17, 1.31067438509808e+17, 1.31067438514183e+17, 1.31067438518558e+17, 1.310674385226205e+17, 1.31067438526683e+17, 1.310674385312143e+17, 1.310674385352767e+17, 1.310674385394954e+17, 1.31067438543558e+17, 1.310674385476205e+17, 1.310674385516829e+17, 1.310674385559017e+17, 1.310674385599643e+17, 1.310674385640268e+17, 1.310674385680892e+17, 1.31067438572308e+17, 1.31067438576683e+17, 1.31067438581058e+17, 1.310674385855892e+17, 1.310674385896517e+17, 1.310674385937143e+17, 1.310674385984017e+17, 1.310674386024643e+17, 1.310674386065267e+17, 1.310674386107456e+17, 1.310674386149642e+17, 1.310674386193393e+17, 1.310674386234017e+17, 1.310674386277768e+17, 1.310674386319955e+17, 1.31067438636058e+17, 1.310674386405893e+17, 1.310674386448081e+17, 1.310674386488704e+17, 1.31067438652933e+17, 1.310674386576205e+17, 1.31067438662308e+17, 1.310674386668393e+17, 1.310674386709018e+17, 1.310674386749642e+17, 1.310674386790268e+17, 1.310674386830893e+17, 1.310674386871517e+17, 1.310674386912142e+17, 1.31067438695433e+17, 1.31067438699808e+17, 1.310674387038705e+17, 1.310674387079331e+17, 1.310674387124643e+17, 1.310674387165267e+17, 1.310674387207456e+17, 1.310674387251205e+17, 1.310674387293393e+17, 1.31067438733558e+17, 1.310674387377768e+17, 1.31067438742308e+17, 1.310674387469955e+17, 1.31067438751058e+17, 1.310674387551205e+17, 1.310674387593393e+17, 1.310674387632456e+17, 1.310674387673079e+17, 1.310674387713705e+17, 1.310674387754331e+17, 1.310674387794954e+17, 1.31067438783558e+17, 1.310674387876205e+17, 1.310674387918394e+17, 1.310674387959017e+17, 1.310674387999643e+17, 1.310674388044955e+17, 1.31067438808558e+17, 1.310674388126205e+17, 1.310674388168393e+17, 1.310674388209018e+17, 1.310674388251205e+17, 1.310674388293393e+17, 1.31067438833558e+17, 1.310674388379331e+17, 1.310674388419955e+17, 1.310674388463704e+17, 1.31067438850433e+17, 1.310674388544955e+17, 1.310674388587142e+17, 1.310674388627767e+17, 1.310674388669955e+17, 1.310674388713705e+17, 1.310674388757455e+17, 1.31067438879808e+17, 1.310674388838705e+17, 1.310674388880892e+17, 1.310674388924643e+17, 1.310674388965267e+17, 1.31067438900433e+17, 1.310674389044955e+17, 1.310674389085581e+17, 1.310674389126205e+17, 1.310674389168393e+17, 1.310674389207455e+17, 1.310674389251205e+17, 1.31067438929183e+17, 1.310674389332454e+17, 1.310674389380892e+17, 1.31067438942308e+17, 1.310674389465267e+17, 1.310674389507455e+17, 1.310674389549642e+17, 1.310674389590267e+17, 1.310674389634017e+17, 1.310674389677768e+17, 1.310674389718392e+17, 1.310674389759017e+17, 1.310674389799642e+17, 1.31067438984183e+17, 1.310674389884017e+17, 1.310674389924643e+17, 1.310674389968392e+17, 1.31067439001058e+17, 1.31067439005433e+17, 1.310674390096517e+17, 1.310674390140268e+17, 1.310674390182455e+17, 1.31067439022308e+17, 1.310674390263706e+17, 1.310674390302767e+17, 1.310674390343393e+17, 1.310674390388704e+17, 1.310674390427768e+17, 1.310674390468393e+17, 1.310674390512143e+17, 1.310674390552767e+17, 1.310674390593393e+17, 1.31067439063558e+17, 1.310674390676205e+17, 1.310674390715268e+17, 1.310674390755892e+17, 1.310674390796517e+17, 1.310674390837142e+17, 1.310674390877768e+17, 1.310674390919955e+17, 1.31067439096058e+17, 1.310674391001204e+17, 1.31067439104183e+17, 1.310674391084018e+17, 1.310674391124643e+17, 1.310674391165267e+17, 1.310674391207455e+17, 1.310674391248081e+17, 1.310674391288705e+17, 1.31067439132933e+17, 1.310674391369956e+17, 1.31067439141058e+17, 1.310674391455892e+17, 1.310674391496517e+17, 1.310674391537142e+17, 1.310674391577768e+17, 1.310674391618394e+17, 1.310674391662143e+17, 1.310674391702769e+17, 1.310674391743392e+17, 1.310674391784017e+17, 1.310674391826205e+17, 1.310674391869955e+17, 1.31067439191058e+17, 1.310674391951205e+17, 1.31067439199808e+17, 1.310674392038705e+17, 1.310674392080893e+17, 1.310674392126204e+17, 1.31067439216683e+17, 1.310674392207455e+17, 1.310674392248079e+17, 1.310674392288705e+17, 1.310674392327768e+17, 1.310674392368393e+17, 1.310674392409018e+17, 1.310674392451205e+17, 1.310674392494954e+17, 1.31067439253558e+17, 1.310674392577768e+17, 1.310674392618392e+17, 1.310674392659017e+17, 1.310674392699643e+17, 1.310674392740268e+17, 1.310674392779331e+17, 1.310674392819955e+17, 1.31067439286058e+17, 1.31067439290433e+17, 1.310674392944955e+17, 1.31067439298558e+17, 1.310674393027768e+17, 1.310674393068392e+17, 1.310674393109018e+17, 1.310674393149642e+17, 1.310674393190268e+17, 1.310674393230893e+17, 1.310674393271517e+17, 1.310674393312143e+17, 1.310674393352767e+17, 1.310674393393393e+17, 1.310674393434019e+17, 1.310674393476205e+17, 1.310674393516829e+17, 1.310674393557455e+17, 1.310674393596517e+17, 1.310674393637143e+17, 1.310674393677768e+17, 1.31067439372308e+17, 1.310674393765267e+17, 1.310674393809016e+17, 1.310674393851205e+17, 1.310674393896518e+17, 1.310674393937142e+17, 1.310674393977768e+17, 1.310674394021517e+17, 1.310674394062143e+17, 1.310674394102767e+17},
			             {1.310674180084018e+17, 1.310674180376205e+17},
			             {1.31067417557308e+17, 1.310674175774642e+17},
			             {1.310674183543392e+17, 1.310674183676205e+17},
			             {1.310674184707456e+17, 1.310674184869955e+17},
			             {1.310674305199643e+17, 1.310674305362141e+17},
			             {1.310674306415268e+17, 1.310674306459018e+17, 1.310674306499643e+17, 1.31067430654183e+17, 1.310674306584018e+17, 1.31067430662933e+17, 1.310674306671517e+17, 1.310674306712143e+17, 1.310674306752768e+17, 1.31067430679808e+17, 1.310674306838705e+17, 1.310674306879329e+17, 1.310674306921518e+17, 1.310674306962143e+17, 1.310674307002767e+17, 1.310674307048081e+17, 1.310674307088705e+17, 1.31067430712933e+17, 1.310674307169956e+17, 1.31067430721058e+17, 1.310674307259018e+17, 1.310674307302767e+17, 1.310674307343392e+17},
			             {1.310674275344955e+17, 1.310674275480893e+17},
			             {1.310674275302767e+17, 1.310674275480893e+17},
			             {1.310674276437143e+17, 1.310674276685581e+17},
			             {1.31067427949183e+17, 1.310674279699643e+17},
			             {1.31067422176683e+17, 1.310674221807456e+17, 1.310674221848079e+17, 1.310674221890267e+17, 1.310674221971517e+17, 1.310674222012142e+17, 1.31067422206058e+17, 1.310674222101204e+17},
			             {1.310674231143392e+17, 1.310674231309018e+17},
			             {1.310674196838706e+17, 1.310674197084017e+17},
			             {1.310674242009018e+17, 1.310674242140268e+17},
			             {1.310674257349642e+17, 1.310674257469956e+17},
			             {1.310674260618392e+17, 1.310674260743393e+17},
			             {1.310674310044955e+17, 1.310674310219955e+17},
			             {1.310674313924643e+17, 1.310674314132454e+17},
			             {1.31067431426683e+17, 1.310674314515268e+17},
			             {1.310674316476205e+17, 1.310674316601204e+17},
			             {1.310674316857455e+17, 1.310674317024643e+17},
			             {1.310674248162143e+17, 1.310674248284018e+17},
			             {1.310674322724643e+17, 1.31067432289183e+17, 1.310674322938706e+17},
			             {1.310674323319954e+17, 1.310674323571517e+17},
			             {1.310674325077768e+17, 1.310674325321517e+17},
			             {1.310674329571517e+17, 1.310674329779331e+17};
			mask_depths = {{15.0, 15.0, 52.6, 52.6}, {15.0, 52.5}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.6}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.7}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.8}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 52.9}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.0}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.1}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.2}, {15.0, 53.2}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.6}, {15.0, 53.5}, {15.0, 53.6}, {15.0, 53.7}, {15.0, 53.7}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.3}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.5}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.5}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.4}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.5}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.7}, {15.0, 53.6}, {15.0, 53.7}, {15.0, 53.7}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.7}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.6}, {15.0, 53.7}, {15.0, 53.7}, {15.0, 53.7}, {15.0, 53.7}, {15.0, 53.7}, {15.0, 53.7}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.8}, {15.0, 53.8}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.3}, {15.0, 54.2}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.4}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.7}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.8}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.8}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.0}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.1}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.3}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.3}, {15.0, 55.2}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.5}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.9}, {15.0, 55.8}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.7}, {15.0, 56.8}, {15.0, 56.7}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.8}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.8}, {15.0, 56.9}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.1}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.3}, {15.0, 57.2}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.5}, {15.0, 57.6}, {15.0, 57.5}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.7}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.8}, {15.0, 57.9}, {15.0, 57.8}, {15.0, 57.9}, {15.0, 57.8}, {15.0, 57.9}, {15.0, 58.0}, {15.0, 58.0}, {15.0, 58.1}, {15.0, 58.0}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.0}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.0}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.0}, {15.0, 58.0}, {15.0, 58.0}, {15.0, 58.0}, {15.0, 58.1}, {15.0, 58.0}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.1}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.1}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.5}, {15.0, 58.4}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.4}, {15.0, 58.5}, {15.0, 58.4}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.7}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.7}, {15.0, 58.7}, {15.0, 58.7}, {15.0, 58.8}, {15.0, 58.7}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.1}, {15.0, 59.2}, {15.0, 59.1}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.4}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.1}, {15.0, 59.2}, {15.0, 59.1}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.4}, {15.0, 59.4}, {15.0, 59.4}, {15.0, 59.4}, {15.0, 59.4}, {15.0, 59.5}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.5}, {15.0, 59.6}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.4}, {15.0, 59.5}, {15.0, 59.4}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.7}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.9}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.7}, {15.0, 59.8}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.2}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.2}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.2}, {15.0, 60.2}, {15.0, 60.2}, {15.0, 60.2}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.3}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.5}, {15.0, 60.6}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.6}, {15.0, 60.5}, {15.0, 60.6}, {15.0, 60.5}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.5}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.2}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.2}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.1}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 61.0}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.7}, {15.0, 61.7}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.7}, {15.0, 61.7}, {15.0, 61.7}, {15.0, 61.7}, {15.0, 61.6}, {15.0, 61.6}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.3}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.4}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 61.5}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 15.0, 60.7, 60.7}}, {{15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.9}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.8}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.7}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.6}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.4}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.5}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.4}, {15.0, 60.3}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.4}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.2}, {15.0, 60.2}, {15.0, 60.2}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.2}, {15.0, 60.2}, {15.0, 60.2}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.2}, {15.0, 60.3}, {15.0, 60.2}, {15.0, 60.2}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.1}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.1}, {15.0, 60.0}, {15.0, 60.1}, {15.0, 60.1}, {15.0, 60.0}, {15.0, 60.1}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.7}, {15.0, 59.6}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.8}, {15.0, 59.8}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 60.0}, {15.0, 59.9}, {15.0, 59.9}, {15.0, 59.8}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.4}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.7}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.6}, {15.0, 59.5}, {15.0, 59.4}, {15.0, 59.4}, {15.0, 59.4}, {15.0, 59.3}, {15.0, 59.4}, {15.0, 59.4}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.4}, {15.0, 59.4}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.5}, {15.0, 59.4}, {15.0, 59.3}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.3}, {15.0, 59.2}, {15.0, 59.3}, {15.0, 59.3}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.2}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.0}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.9}, {15.0, 59.0}, {15.0, 58.9}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.1}, {15.0, 59.1}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 59.0}, {15.0, 58.9}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.7}, {15.0, 58.7}, {15.0, 58.7}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.7}, {15.0, 58.7}, {15.0, 58.7}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.8}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.9}, {15.0, 58.8}, {15.0, 58.7}, {15.0, 58.7}, {15.0, 58.6}, {15.0, 58.6}, {15.0, 58.5}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.4}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.5}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.4}, {15.0, 58.3}, {15.0, 58.4}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.2}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.2}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.2}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.3}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.0}, {15.0, 58.0}, {15.0, 58.0}, {15.0, 58.0}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.2}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.1}, {15.0, 58.0}, {15.0, 58.0}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.9}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.9}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.9}, {15.0, 57.8}, {15.0, 57.8}, {15.0, 57.9}, {15.0, 57.8}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.7}, {15.0, 57.7}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.6}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.6}, {15.0, 57.5}, {15.0, 57.6}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.5}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.4}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.3}, {15.0, 57.2}, {15.0, 57.2}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.1}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 57.0}, {15.0, 56.9}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.7}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.7}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.9}, {15.0, 56.8}, {15.0, 56.8}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.6}, {15.0, 56.7}, {15.0, 56.6}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.7}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.6}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.4}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.5}, {15.0, 56.4}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.3}, {15.0, 56.4}, {15.0, 56.3}, {15.0, 56.4}, {15.0, 56.4}, {15.0, 56.3}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.3}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.2}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 55.9}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.7}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 56.0}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.1}, {15.0, 56.2}, {15.0, 56.1}, {15.0, 56.2}, {15.0, 56.1}, {15.0, 56.2}, {15.0, 56.1}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 56.0}, {15.0, 55.9}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 56.0}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.8}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.9}, {15.0, 55.8}, {15.0, 55.9}, {15.0, 55.8}, {15.0, 55.8}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.7}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.7}, {15.0, 55.6}, {15.0, 55.7}, {15.0, 55.6}, {15.0, 55.7}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.7}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.6}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.5}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.2}, {15.0, 55.3}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.4}, {15.0, 55.3}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.3}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.0}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.2}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.0}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.2}, {15.0, 55.1}, {15.0, 55.1}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 55.0}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.8}, {15.0, 54.9}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.9}, {15.0, 54.8}, {15.0, 54.8}, {15.0, 54.7}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.7}, {15.0, 54.8}, {15.0, 54.7}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.6}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.5}, {15.0, 54.5}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.4}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.3}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.3}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.3}, {15.0, 54.2}, {15.0, 54.3}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 53.9}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.0}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.2}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 54.1}, {15.0, 15.0, 54.1, 54.1}}, {{45.2, 50.0}, {45.2, 50.0}}, {{32.9, 35.8}, {32.9, 35.8}}, {{40.3, 44.2}, {40.3, 44.2}}, {{49.1, 51.7}, {49.1, 51.7}}, {{47.4, 52.1}, {47.4, 52.1}}, {{49.1, 54.9}, {55.0, 55.3}, {55.4, 55.7}, {55.8, 56.0}, {56.1, 56.3}, {56.4, 56.7}, {56.8, 57.1}, {57.2, 57.3}, {57.4, 57.5}, {57.6, 57.8}, {49.1, 49.4, 57.9, 58.0}, {49.5, 50.1, 58.1, 58.4}, {50.2, 50.6}, {50.7, 51.1, 58.6, 58.7}, {51.2, 51.8, 58.8, 59.0}, {51.9, 52.1, 59.1, 59.2}, {52.2, 52.6, 59.3, 59.4}, {52.7, 52.9}, {53.0, 53.4}, {53.5, 54.4}, {54.5, 54.8}, {54.9, 55.2}, {55.3, 59.4}}, {{41.2, 48.3}, {41.2, 48.3}}, {{51.7, 57.8}, {51.7, 57.8}}, {{48.1, 55.2}, {48.1, 55.2}}, {{49.2, 53.3}, {49.2, 53.3}}, {{51.6, 54.5}, {54.4}, {54.4}, {54.5}, {54.5}, {54.6}, {54.5}, {51.6, 54.5}}, {{45.7, 52.9}, {45.7, 52.9}}, {{47.8, 50.7}, {47.8, 50.7}}, {{49.9, 52.8}, {49.9, 52.8}}, {{52.3, 56.0}, {52.3, 56.0}}, {{46.4, 52.0}, {46.4, 52.0}}, {{52.2, 55.9}, {52.2, 55.9}}, {{55.9, 58.1}, {55.9, 58.1}}, {{50.8, 55.7}, {50.8, 55.7}}, {{49.7, 53.6}, {49.7, 53.6}}, {{58.5, 60.3}, {58.5, 60.3}}, {{55.5, 58.8}, {55.5, 58.8}}, {{59.4, 61.4}, {61.4}, {59.4, 61.3}}, {{53.6, 58.7}, {53.6, 58.7}}, {{48.3, 58.3}, {48.3, 58.3}}, {{51.9, 55.8}, {51.9, 55.8}};
		}
	}
}
