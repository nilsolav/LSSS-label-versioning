netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200729T093456";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 4;
			channels = 6;
			categories = 24;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0, 23.5, 38.8,  2.2;
			max_depth =  58.5, 25.8, 43.2,  3.1;
			start_time = 131381358480950784, 131381364866107008, 131381378687825792, 131381380969232000;
			end_time = 131381380969232000, 131381364884700800, 131381378708606976, 131381380969232000;
			region_id = 1, 2, 3, 4;
			region_name = "Layer1","Layer1","Layer2","Layer3";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "";
			region_category_names = "0", "0", "0", "0", "0", "0", "1", "1", "1", "1", "1", "1", "27", "27", "27", "27", "27", "27", "5027", "5027", "5027", "5027", "5027", "5027";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24;
			region_type = analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "333";
			region_channels = 63, 63, 63, 63;
			mask_times = {1.313813584809508e+17, 1.31381358488607e+17, 1.313813584926694e+17, 1.313813584950132e+17, 1.313813585059507e+17, 1.313813585109508e+17, 1.313813585165757e+17, 1.313813585240758e+17, 1.313813585320444e+17, 1.313813585378258e+17, 1.313813585462632e+17, 1.313813585511069e+17, 1.313813585570445e+17, 1.313813585645445e+17, 1.313813585706382e+17, 1.313813585776695e+17, 1.313813585851694e+17, 1.31381358590482e+17, 1.313813585928257e+17, 1.313813586043882e+17, 1.313813586068882e+17, 1.313813586178257e+17, 1.313813586207945e+17, 1.313813586231383e+17, 1.313813586342319e+17, 1.313813586372008e+17, 1.313813586490758e+17, 1.313813586526696e+17, 1.313813586584507e+17, 1.313813586654821e+17, 1.313813586718883e+17, 1.31381358678607e+17, 1.313813586850132e+17, 1.313813586907945e+17, 1.313813586965757e+17, 1.313813587042319e+17, 1.313813587090757e+17, 1.313813587159507e+17, 1.313813587232945e+17, 1.313813587306382e+17, 1.313813587362632e+17, 1.313813587437632e+17, 1.313813587512632e+17, 1.313813587587633e+17, 1.313813587653257e+17, 1.313813587676695e+17, 1.313813587734508e+17, 1.313813587803258e+17, 1.31381358786732e+17, 1.31381358793607e+17, 1.313813587997007e+17, 1.313813588064196e+17, 1.313813588131383e+17, 1.31381358819857e+17, 1.313813588264196e+17, 1.313813588289196e+17, 1.313813588406382e+17, 1.31381358842982e+17, 1.313813588500132e+17, 1.313813588603256e+17, 1.313813588634508e+17, 1.313813588706382e+17, 1.31381358877982e+17, 1.313813588887633e+17, 1.31381358892982e+17, 1.313813589012634e+17, 1.313813589093883e+17, 1.313813589142321e+17, 1.313813589173569e+17, 1.31381358922357e+17, 1.313813589331382e+17, 1.313813589400133e+17, 1.313813589473571e+17, 1.313813589543882e+17, 1.313813589606382e+17, 1.313813589676695e+17, 1.313813589734508e+17, 1.313813589803258e+17, 1.313813589862633e+17, 1.313813589934508e+17, 1.31381359000482e+17, 1.313813590087633e+17, 1.31381359018607e+17, 1.313813590222007e+17, 1.313813590289196e+17, 1.313813590353257e+17, 1.313813590434508e+17, 1.313813590504819e+17, 1.313813590579821e+17, 1.313813590678257e+17, 1.313813590728257e+17, 1.31381359079857e+17, 1.313813590851695e+17, 1.313813590931383e+17, 1.31381359099232e+17, 1.313813591062632e+17, 1.31381359112357e+17, 1.313813591201695e+17, 1.313813591225133e+17, 1.313813591340758e+17, 1.313813591364196e+17, 1.313813591443882e+17, 1.313813591512632e+17, 1.31381359159232e+17, 1.313813591659507e+17, 1.313813591725133e+17, 1.313813591789196e+17, 1.313813591847007e+17, 1.313813591907944e+17, 1.313813591981382e+17, 1.313813592100132e+17, 1.313813592132945e+17, 1.313813592207945e+17, 1.313813592262633e+17, 1.313813592343882e+17, 1.313813592414195e+17, 1.313813592493883e+17, 1.313813592570445e+17, 1.313813592672008e+17, 1.313813592756383e+17, 1.313813592807945e+17, 1.313813592882945e+17, 1.313813592943884e+17, 1.313813593009508e+17, 1.313813593082945e+17, 1.31381359315482e+17, 1.313813593243882e+17, 1.313813593331383e+17, 1.313813593418883e+17, 1.313813593456383e+17, 1.31381359347982e+17, 1.31381359359857e+17, 1.313813593622007e+17, 1.313813593731383e+17, 1.313813593787633e+17, 1.313813593875132e+17, 1.313813593972008e+17, 1.313813594050132e+17, 1.313813594137632e+17, 1.313813594197007e+17, 1.313813594273571e+17, 1.31381359436107e+17, 1.313813594443884e+17, 1.313813594490757e+17, 1.313813594559507e+17, 1.313813594612632e+17, 1.313813594686071e+17, 1.313813594725133e+17, 1.313813594806382e+17, 1.313813594875132e+17, 1.313813594939195e+17, 1.313813595003258e+17, 1.313813595075133e+17, 1.313813595134508e+17, 1.313813595207945e+17, 1.31381359527982e+17, 1.313813595348571e+17, 1.31381359542357e+17, 1.313813595481382e+17, 1.313813595543884e+17, 1.313813595614195e+17, 1.31381359566107e+17, 1.313813595750132e+17, 1.313813595773571e+17, 1.313813595897007e+17, 1.313813595962633e+17, 1.313813596011071e+17, 1.313813596084508e+17, 1.313813596157946e+17, 1.313813596239195e+17, 1.31381359632982e+17, 1.313813596378257e+17, 1.313813596442321e+17, 1.313813596500132e+17, 1.313813596568883e+17, 1.313813596642321e+17, 1.313813596712632e+17, 1.313813596772008e+17, 1.313813596851695e+17, 1.313813596925133e+17, 1.313813597014195e+17, 1.313813597062633e+17, 1.313813597120444e+17, 1.313813597189196e+17, 1.313813597262633e+17, 1.313813597332945e+17, 1.313813597397007e+17, 1.313813597468883e+17, 1.313813597542321e+17, 1.313813597614195e+17, 1.313813597693883e+17, 1.31381359778607e+17, 1.313813597809508e+17, 1.31381359784857e+17, 1.313813597942321e+17, 1.313813598001695e+17, 1.313813598072008e+17, 1.313813598132945e+17, 1.31381359820482e+17, 1.313813598278258e+17, 1.31381359836107e+17, 1.31381359842357e+17, 1.31381359846732e+17, 1.313813598490757e+17, 1.313813598611071e+17, 1.31381359866107e+17, 1.31381359872357e+17, 1.313813598789194e+17, 1.313813598850132e+17, 1.313813598918883e+17, 1.313813598995444e+17, 1.313813599059507e+17, 1.31381359909857e+17, 1.313813599170445e+17, 1.313813599239195e+17, 1.313813599309508e+17, 1.313813599332945e+17, 1.313813599457944e+17, 1.31381359952982e+17, 1.313813599603258e+17, 1.313813599670445e+17, 1.313813599745445e+17, 1.313813599768882e+17, 1.31381359989232e+17, 1.313813599922007e+17, 1.31381359999232e+17, 1.313813600034508e+17, 1.313813600109507e+17, 1.31381360019232e+17, 1.31381360027982e+17, 1.313813600328257e+17, 1.313813600397007e+17, 1.313813600465757e+17, 1.313813600532945e+17, 1.313813600557944e+17, 1.31381360065482e+17, 1.313813600718883e+17, 1.313813600800133e+17, 1.313813600853257e+17, 1.313813600920445e+17, 1.313813600979821e+17, 1.313813601068882e+17, 1.313813601129819e+17, 1.313813601190757e+17, 1.31381360126107e+17, 1.313813601332945e+17, 1.313813601400133e+17, 1.313813601476695e+17, 1.313813601542319e+17, 1.313813601634508e+17, 1.31381360166732e+17, 1.313813601740758e+17, 1.313813601812632e+17, 1.313813601887633e+17, 1.313813601976695e+17, 1.313813602014195e+17, 1.313813602081382e+17, 1.313813602150132e+17, 1.313813602232945e+17, 1.313813602306383e+17, 1.313813602375132e+17, 1.313813602465757e+17, 1.31381360253607e+17, 1.313813602582945e+17, 1.313813602678257e+17, 1.313813602717321e+17, 1.313813602779821e+17, 1.313813602831382e+17, 1.31381360290482e+17, 1.313813602976695e+17, 1.313813603037632e+17, 1.313813603112634e+17, 1.313813603175132e+17, 1.313813603247008e+17, 1.313813603342321e+17, 1.313813603414194e+17, 1.313813603439195e+17, 1.313813603504819e+17, 1.313813603562633e+17, 1.313813603643882e+17, 1.313813603726696e+17, 1.313813603775132e+17, 1.313813603853258e+17, 1.31381360392982e+17, 1.313813604001695e+17, 1.313813604072008e+17, 1.313813604143882e+17, 1.313813604226694e+17, 1.313813604301695e+17, 1.31381360438607e+17, 1.313813604442321e+17, 1.313813604465757e+17, 1.31381360459232e+17, 1.31381360462982e+17, 1.313813604718883e+17, 1.31381360479232e+17, 1.313813604873571e+17, 1.313813604920444e+17, 1.313813605039195e+17, 1.313813605082944e+17, 1.313813605159508e+17, 1.31381360521732e+17, 1.313813605240758e+17, 1.313813605362633e+17, 1.313813605401695e+17, 1.31381360548607e+17, 1.31381360556732e+17, 1.313813605701696e+17, 1.313813605725133e+17, 1.313813605750132e+17, 1.31381360584857e+17, 1.313813605873569e+17, 1.313813605987633e+17, 1.313813606057946e+17, 1.313813606120445e+17, 1.313813606195444e+17, 1.313813606268882e+17, 1.313813606340756e+17, 1.313813606414195e+17, 1.313813606481382e+17, 1.313813606506382e+17, 1.313813606565757e+17, 1.313813606657944e+17, 1.313813606728257e+17, 1.313813606803256e+17, 1.313813606875132e+17, 1.313813607001695e+17, 1.313813607025133e+17, 1.31381360709857e+17, 1.31381360716107e+17, 1.31381360723607e+17, 1.313813607309508e+17, 1.313813607381382e+17, 1.313813607500133e+17, 1.313813607540758e+17, 1.313813607603258e+17, 1.313813607664196e+17, 1.313813607748571e+17, 1.31381360782357e+17, 1.313813607881382e+17, 1.313813607962633e+17, 1.313813607987633e+17, 1.31381360809857e+17, 1.313813608140756e+17, 1.313813608218883e+17, 1.313813608304819e+17, 1.313813608356383e+17, 1.31381360841732e+17, 1.313813608440758e+17, 1.313813608573571e+17, 1.313813608650132e+17, 1.313813608704819e+17, 1.313813608728257e+17, 1.313813608851694e+17, 1.313813608914195e+17, 1.313813608990757e+17, 1.313813609072008e+17, 1.313813609145445e+17, 1.313813609220445e+17, 1.313813609295444e+17, 1.313813609320445e+17, 1.313813609447007e+17, 1.313813609511069e+17, 1.313813609584507e+17, 1.313813609656383e+17, 1.313813609742319e+17, 1.31381360982982e+17, 1.313813609881382e+17, 1.31381360990482e+17, 1.313813610029819e+17, 1.313813610056383e+17, 1.313813610120444e+17, 1.313813610193882e+17, 1.31381361026107e+17, 1.31381361032982e+17, 1.31381361039857e+17, 1.313813610470445e+17, 1.313813610493883e+17, 1.313813610615758e+17, 1.313813610709508e+17, 1.313813610753257e+17, 1.313813610778258e+17, 1.313813610893883e+17, 1.313813610976695e+17, 1.313813611020444e+17, 1.313813611043882e+17, 1.31381361116732e+17, 1.31381361120482e+17, 1.313813611257946e+17, 1.313813611309508e+17, 1.31381361136732e+17, 1.313813611451694e+17, 1.313813611525133e+17, 1.313813611595444e+17, 1.313813611664195e+17, 1.313813611747008e+17, 1.313813611789196e+17, 1.313813611857944e+17, 1.313813611922008e+17, 1.313813612004819e+17, 1.313813612075132e+17, 1.313813612109508e+17, 1.313813612218883e+17, 1.313813612303258e+17, 1.313813612364196e+17, 1.313813612422007e+17, 1.313813612501695e+17, 1.31381361256732e+17, 1.313813612634508e+17, 1.31381361269857e+17, 1.313813612773571e+17, 1.313813612857946e+17, 1.31381361292357e+17, 1.313813612993883e+17, 1.313813613075133e+17, 1.313813613178258e+17, 1.313813613232945e+17, 1.313813613303258e+17, 1.313813613328257e+17, 1.31381361344857e+17, 1.313813613553257e+17, 1.313813613579821e+17, 1.313813613640758e+17, 1.313813613681382e+17, 1.31381361374857e+17, 1.313813613815758e+17, 1.313813613890757e+17, 1.313813613965757e+17, 1.313813614037633e+17, 1.313813614101696e+17, 1.313813614182945e+17, 1.313813614242321e+17, 1.313813614322007e+17, 1.313813614448571e+17, 1.313813614473571e+17, 1.313813614556383e+17, 1.313813614614195e+17, 1.31381361469232e+17, 1.31381361476732e+17, 1.313813614840756e+17, 1.313813614953257e+17, 1.313813614997007e+17, 1.313813615078257e+17, 1.313813615172008e+17, 1.313813615228257e+17, 1.313813615312632e+17, 1.313813615415757e+17, 1.313813615468883e+17, 1.31381361549232e+17, 1.31381361561732e+17, 1.313813615693883e+17, 1.31381361571732e+17, 1.313813615845445e+17, 1.313813615928257e+17, 1.313813616000133e+17, 1.313813616103258e+17, 1.313813616140758e+17, 1.31381361621732e+17, 1.313813616290757e+17, 1.313813616364195e+17, 1.313813616439195e+17, 1.313813616506382e+17, 1.313813616576695e+17, 1.313813616650132e+17, 1.313813616722008e+17, 1.313813616790757e+17, 1.313813616851695e+17, 1.313813616937632e+17, 1.313813617003258e+17, 1.313813617084508e+17, 1.313813617151695e+17, 1.31381361722982e+17, 1.313813617290757e+17, 1.313813617314195e+17, 1.313813617439195e+17, 1.313813617490757e+17, 1.31381361756107e+17, 1.313813617634508e+17, 1.313813617734508e+17, 1.313813617757944e+17, 1.31381361786107e+17, 1.313813617900133e+17, 1.313813617976695e+17, 1.313813618064196e+17, 1.31381361810482e+17, 1.313813618197007e+17, 1.31381361824857e+17, 1.313813618322007e+17, 1.313813618395444e+17, 1.313813618467319e+17, 1.31381361852357e+17, 1.313813618547007e+17, 1.313813618675132e+17, 1.313813618756383e+17, 1.31381361882982e+17, 1.313813618912632e+17, 1.313813618997007e+17, 1.313813619070445e+17, 1.313813619126696e+17, 1.313813619225133e+17, 1.313813619287633e+17, 1.313813619362633e+17, 1.313813619437632e+17, 1.313813619520445e+17, 1.313813619604819e+17, 1.313813619679821e+17, 1.313813619775132e+17, 1.313813619828257e+17, 1.313813619906382e+17, 1.31381361998607e+17, 1.313813620032945e+17, 1.313813620132945e+17, 1.313813620195446e+17, 1.31381362026732e+17, 1.313813620340758e+17, 1.313813620422008e+17, 1.313813620473569e+17, 1.313813620545445e+17, 1.313813620612632e+17, 1.313813620695444e+17, 1.313813620768882e+17, 1.313813620842319e+17, 1.313813620901695e+17, 1.313813620978258e+17, 1.31381362106107e+17, 1.313813621109508e+17, 1.313813621187633e+17, 1.313813621265757e+17, 1.313813621328257e+17, 1.31381362136732e+17, 1.313813621437632e+17, 1.31381362151732e+17, 1.313813621576695e+17, 1.313813621650132e+17, 1.313813621722007e+17, 1.31381362180482e+17, 1.313813621870445e+17, 1.313813621943882e+17, 1.313813622007945e+17, 1.313813622081382e+17, 1.313813622156383e+17, 1.31381362222982e+17, 1.313813622314195e+17, 1.313813622387633e+17, 1.313813622470445e+17, 1.313813622553258e+17, 1.313813622626696e+17, 1.31381362269857e+17, 1.313813622800132e+17, 1.313813622857946e+17, 1.313813622920444e+17, 1.313813622993883e+17, 1.31381362304857e+17, 1.31381362314857e+17, 1.313813623220445e+17, 1.31381362330482e+17, 1.313813623378258e+17, 1.313813623465757e+17, 1.313813623528257e+17, 1.31381362360482e+17, 1.313813623675132e+17, 1.31381362369857e+17, 1.313813623822008e+17, 1.313813623893883e+17, 1.313813624006382e+17, 1.313813624040758e+17, 1.313813624064195e+17, 1.313813624151695e+17, 1.313813624215757e+17, 1.313813624351695e+17, 1.313813624375133e+17, 1.313813624451694e+17, 1.31381362450482e+17, 1.313813624587633e+17, 1.31381362466107e+17, 1.313813624732945e+17, 1.313813624837633e+17, 1.31381362486732e+17, 1.31381362489232e+17, 1.313813624995446e+17, 1.31381362505482e+17, 1.313813625128257e+17, 1.313813625200132e+17, 1.313813625265757e+17, 1.313813625337632e+17, 1.313813625412632e+17, 1.313813625484507e+17, 1.313813625557944e+17, 1.313813625618883e+17, 1.313813625642319e+17, 1.313813625773571e+17, 1.313813625825133e+17, 1.313813625907945e+17, 1.313813625931383e+17, 1.313813626051695e+17, 1.313813626089196e+17, 1.313813626128257e+17, 1.313813626231383e+17, 1.313813626312632e+17, 1.313813626384507e+17, 1.313813626462633e+17, 1.313813626500132e+17, 1.313813626573571e+17, 1.313813626648571e+17, 1.313813626712632e+17, 1.313813626803256e+17, 1.31381362685482e+17, 1.31381362692982e+17, 1.313813627022007e+17, 1.313813627075132e+17, 1.31381362709857e+17, 1.313813627218883e+17, 1.313813627242321e+17, 1.313813627286071e+17, 1.313813627393883e+17, 1.313813627465757e+17, 1.313813627537632e+17, 1.313813627600133e+17, 1.313813627665756e+17, 1.313813627739195e+17, 1.313813627809508e+17, 1.313813627881382e+17, 1.313813627947008e+17, 1.313813628012632e+17, 1.313813628103258e+17, 1.313813628153258e+17, 1.313813628176695e+17, 1.31381362829857e+17, 1.313813628343882e+17, 1.313813628414195e+17, 1.313813628509508e+17, 1.313813628540756e+17, 1.313813628609508e+17, 1.313813628657946e+17, 1.313813628745445e+17, 1.313813628784507e+17, 1.31381362885482e+17, 1.313813628926696e+17, 1.313813628950132e+17, 1.313813629078258e+17, 1.313813629103258e+17, 1.313813629164196e+17, 1.313813629222007e+17, 1.313813629293883e+17, 1.313813629365757e+17, 1.313813629428257e+17, 1.31381362949857e+17, 1.313813629522007e+17, 1.313813629643882e+17, 1.31381362966732e+17, 1.313813629745445e+17, 1.313813629811069e+17, 1.313813629893883e+17, 1.313813629950132e+17, 1.313813630022007e+17, 1.31381363009232e+17, 1.313813630164196e+17, 1.313813630236069e+17, 1.313813630306382e+17, 1.313813630390757e+17, 1.313813630464195e+17, 1.313813630545445e+17, 1.313813630615757e+17, 1.313813630687633e+17, 1.313813630770445e+17, 1.313813630843882e+17, 1.313813630914195e+17, 1.313813630981382e+17, 1.31381363105482e+17, 1.31381363113607e+17, 1.313813631189194e+17, 1.313813631265757e+17, 1.31381363133607e+17, 1.313813631407945e+17, 1.313813631470446e+17, 1.313813631540756e+17, 1.313813631612632e+17, 1.313813631687631e+17, 1.313813631757946e+17, 1.31381363183607e+17, 1.313813631876695e+17, 1.313813631950132e+17, 1.313813632020444e+17, 1.313813632112632e+17, 1.313813632147008e+17, 1.313813632211071e+17, 1.313813632278258e+17, 1.313813632350132e+17, 1.313813632418883e+17, 1.313813632503258e+17, 1.313813632576695e+17, 1.313813632657944e+17, 1.313813632731382e+17, 1.313813632801696e+17, 1.313813632886071e+17, 1.313813632957944e+17, 1.313813633028257e+17, 1.313813633051695e+17, 1.313813633172008e+17, 1.31381363325482e+17, 1.313813633315757e+17, 1.313813633397007e+17, 1.313813633468883e+17, 1.313813633540756e+17, 1.313813633620445e+17, 1.31381363369232e+17, 1.313813633765757e+17, 1.313813633850132e+17, 1.313813633901696e+17, 1.313813633965757e+17, 1.313813634039195e+17, 1.313813634137633e+17, 1.31381363416732e+17, 1.313813634243882e+17, 1.313813634309508e+17, 1.313813634373571e+17, 1.313813634431383e+17, 1.313813634493883e+17, 1.313813634553257e+17, 1.313813634625133e+17, 1.313813634714195e+17, 1.313813634801695e+17, 1.313813634825133e+17, 1.313813634895444e+17, 1.313813634975132e+17, 1.313813635047007e+17, 1.313813635115758e+17, 1.313813635176695e+17, 1.313813635200133e+17, 1.313813635307944e+17, 1.313813635347008e+17, 1.313813635370445e+17, 1.313813635487633e+17, 1.313813635522008e+17, 1.313813635590757e+17, 1.31381363566732e+17, 1.313813635714195e+17, 1.313813635737632e+17, 1.313813635850132e+17, 1.31381363588607e+17, 1.313813635976695e+17, 1.313813636009508e+17, 1.313813636068883e+17, 1.313813636109507e+17, 1.313813636172008e+17, 1.313813636239195e+17, 1.313813636262632e+17, 1.313813636379821e+17, 1.313813636403258e+17, 1.313813636497007e+17, 1.313813636531383e+17, 1.313813636606382e+17, 1.31381363666107e+17, 1.313813636729819e+17, 1.313813636818883e+17, 1.313813636868882e+17, 1.313813636939195e+17, 1.31381363700482e+17, 1.313813637076695e+17, 1.313813637151695e+17, 1.313813637206383e+17, 1.313813637276695e+17, 1.313813637339195e+17, 1.31381363739857e+17, 1.313813637470445e+17, 1.31381363755482e+17, 1.313813637603258e+17, 1.313813637665757e+17, 1.31381363773607e+17, 1.313813637825133e+17, 1.313813637864195e+17, 1.313813637920444e+17, 1.313813637982945e+17, 1.313813638043882e+17, 1.313813638112632e+17, 1.313813638184508e+17, 1.313813638251695e+17, 1.313813638322007e+17, 1.31381363839232e+17, 1.313813638415757e+17, 1.31381363853607e+17, 1.31381363856107e+17, 1.313813638651695e+17, 1.31381363869232e+17, 1.313813638759507e+17, 1.313813638784508e+17, 1.313813638859508e+17, 1.313813638904819e+17, 1.31381363898607e+17, 1.31381363905482e+17, 1.313813639125133e+17, 1.313813639184507e+17, 1.313813639256383e+17, 1.31381363927982e+17, 1.31381363939232e+17, 1.313813639442321e+17, 1.313813639522007e+17, 1.313813639590757e+17, 1.31381363966732e+17, 1.313813639745445e+17, 1.313813639815757e+17, 1.31381363988607e+17, 1.313813639945445e+17, 1.31381364002357e+17, 1.313813640114195e+17, 1.313813640156383e+17, 1.313813640239195e+17, 1.313813640276695e+17, 1.313813640345445e+17, 1.313813640378258e+17, 1.313813640437633e+17, 1.31381364050482e+17, 1.313813640576695e+17, 1.31381364065482e+17, 1.313813640748571e+17, 1.313813640782945e+17, 1.31381364086732e+17, 1.313813640897007e+17, 1.313813640920444e+17, 1.31381364103607e+17, 1.31381364106107e+17, 1.313813641154821e+17, 1.313813641203258e+17, 1.313813641275132e+17, 1.313813641345445e+17, 1.313813641415758e+17, 1.31381364148607e+17, 1.313813641548571e+17, 1.313813641625133e+17, 1.313813641703258e+17, 1.313813641751695e+17, 1.313813641825133e+17, 1.313813641895444e+17, 1.313813641918883e+17, 1.313813642032945e+17, 1.313813642065757e+17, 1.313813642145445e+17, 1.313813642218883e+17, 1.313813642275132e+17, 1.313813642336069e+17, 1.313813642407945e+17, 1.313813642478258e+17, 1.313813642547008e+17, 1.313813642570445e+17, 1.313813642654821e+17, 1.31381364271732e+17, 1.313813642793883e+17, 1.31381364281732e+17, 1.313813642932945e+17, 1.313813642956381e+17, 1.313813643081382e+17, 1.31381364312982e+17, 1.313813643200132e+17, 1.313813643270445e+17, 1.313813643340758e+17, 1.313813643364195e+17, 1.313813643497007e+17, 1.313813643564195e+17, 1.313813643631382e+17, 1.313813643714195e+17, 1.313813643782944e+17, 1.313813643851695e+17, 1.313813643915757e+17, 1.313813643984508e+17, 1.313813644009508e+17, 1.313813644134508e+17, 1.313813644189196e+17, 1.313813644268882e+17, 1.313813644331383e+17, 1.31381364435482e+17, 1.313813644465757e+17, 1.313813644506382e+17, 1.313813644581382e+17, 1.313813644609507e+17, 1.31381364472357e+17, 1.313813644768883e+17, 1.313813644853258e+17, 1.313813644915758e+17, 1.313813644984508e+17, 1.313813645042321e+17, 1.313813645111069e+17, 1.313813645178257e+17, 1.313813645243884e+17, 1.313813645268882e+17, 1.313813645384508e+17, 1.313813645407945e+17, 1.313813645497007e+17, 1.31381364556732e+17, 1.313813645622007e+17, 1.313813645687633e+17, 1.313813645768882e+17, 1.313813645807945e+17, 1.313813645831383e+17, 1.313813645948571e+17, 1.313813645995446e+17, 1.313813646056383e+17, 1.313813646125133e+17, 1.313813646195444e+17, 1.313813646264196e+17, 1.313813646340756e+17, 1.31381364638607e+17, 1.313813646453257e+17, 1.313813646520444e+17, 1.313813646579821e+17, 1.313813646647008e+17, 1.313813646670445e+17, 1.313813646789196e+17, 1.313813646818883e+17, 1.31381364692982e+17, 1.313813646953257e+17, 1.313813646978257e+17, 1.313813647064195e+17, 1.313813647114195e+17, 1.31381364717982e+17, 1.313813647203256e+17, 1.313813647314195e+17, 1.313813647347008e+17, 1.313813647370445e+17, 1.313813647465757e+17, 1.313813647489194e+17, 1.313813647595444e+17, 1.313813647650132e+17, 1.313813647731382e+17, 1.313813647790757e+17, 1.313813647864195e+17, 1.313813647922008e+17, 1.313813647982945e+17, 1.313813648078257e+17, 1.31381364811732e+17, 1.313813648187633e+17, 1.313813648211069e+17, 1.313813648328257e+17, 1.31381364836732e+17, 1.31381364846107e+17, 1.31381364849232e+17, 1.313813648515757e+17, 1.313813648601695e+17, 1.31381364866107e+17, 1.313813648731383e+17, 1.313813648787633e+17, 1.313813648847008e+17, 1.313813648920445e+17, 1.313813648943884e+17, 1.313813649057946e+17, 1.313813649103258e+17, 1.313813649186071e+17, 1.31381364925482e+17, 1.313813649332945e+17, 1.313813649420444e+17, 1.31381364945482e+17, 1.313813649534508e+17, 1.313813649557946e+17, 1.313813649606382e+17, 1.313813649715758e+17, 1.31381364978607e+17, 1.31381364985482e+17, 1.313813649926696e+17, 1.313813649984507e+17, 1.313813650054821e+17, 1.31381365012357e+17, 1.31381365019232e+17, 1.313813650251695e+17, 1.313813650314195e+17, 1.31381365033607e+17, 1.313813650409508e+17, 1.313813650506382e+17, 1.313813650537632e+17, 1.31381365056107e+17, 1.313813650622007e+17, 1.313813650682944e+17, 1.313813650750132e+17, 1.313813650822008e+17, 1.313813650873571e+17, 1.31381365094857e+17, 1.313813651028257e+17, 1.313813651101695e+17, 1.313813651157944e+17, 1.313813651218883e+17, 1.313813651290757e+17, 1.313813651314195e+17, 1.31381365142982e+17, 1.313813651453257e+17, 1.313813651543884e+17, 1.313813651606382e+17, 1.313813651676695e+17, 1.313813651747007e+17, 1.313813651820444e+17, 1.313813651868882e+17, 1.313813651943884e+17, 1.31381365202357e+17, 1.31381365204857e+17, 1.313813652162633e+17, 1.31381365218607e+17, 1.313813652248571e+17, 1.313813652306382e+17, 1.31381365232982e+17, 1.313813652447008e+17, 1.313813652472008e+17, 1.313813652556383e+17, 1.313813652611071e+17, 1.313813652634508e+17, 1.313813652706382e+17, 1.313813652782945e+17, 1.313813652843882e+17, 1.313813652915758e+17, 1.313813652939195e+17, 1.313813653056383e+17, 1.313813653079821e+17, 1.313813653172008e+17, 1.313813653206382e+17, 1.313813653279821e+17, 1.313813653332945e+17, 1.313813653420445e+17, 1.313813653470445e+17, 1.31381365350482e+17, 1.313813653556383e+17, 1.313813653675133e+17, 1.313813653743882e+17, 1.313813653815758e+17, 1.313813653839196e+17, 1.31381365395482e+17, 1.313813653978258e+17, 1.313813654003258e+17, 1.313813654093883e+17, 1.31381365412357e+17, 1.313813654201695e+17, 1.313813654243882e+17, 1.313813654293883e+17, 1.313813654381382e+17, 1.313813654445445e+17, 1.313813654515757e+17, 1.313813654579821e+17, 1.313813654637632e+17, 1.313813654707945e+17, 1.313813654731383e+17, 1.313813654847008e+17, 1.313813654878258e+17, 1.31381365499857e+17, 1.313813655025133e+17, 1.313813655093882e+17, 1.313813655118883e+17, 1.31381365521732e+17, 1.313813655240756e+17, 1.313813655345445e+17, 1.313813655422007e+17, 1.313813655465757e+17, 1.313813655537632e+17, 1.313813655595444e+17, 1.313813655653257e+17, 1.313813655726694e+17, 1.31381365579857e+17, 1.313813655868883e+17, 1.313813655926694e+17, 1.313813655993883e+17, 1.31381365601732e+17, 1.313813656126694e+17, 1.313813656168882e+17, 1.313813656240758e+17, 1.313813656314195e+17, 1.313813656381382e+17, 1.313813656451695e+17, 1.31381365652357e+17, 1.31381365662982e+17, 1.313813656653258e+17, 1.313813656718883e+17, 1.313813656742321e+17, 1.313813656828257e+17, 1.31381365686732e+17, 1.313813656939195e+17, 1.313813657001695e+17, 1.313813657025133e+17, 1.313813657143884e+17, 1.31381365716732e+17, 1.31381365725482e+17, 1.313813657332945e+17, 1.313813657425133e+17, 1.313813657473571e+17, 1.31381365752982e+17, 1.313813657603256e+17, 1.31381365769232e+17, 1.313813657742321e+17, 1.313813657818883e+17, 1.313813657900133e+17, 1.31381365795482e+17, 1.313813658012634e+17, 1.313813658084507e+17, 1.313813658142321e+17, 1.313813658215757e+17, 1.313813658268883e+17, 1.313813658339195e+17, 1.31381365842982e+17, 1.313813658475133e+17, 1.31381365852357e+17, 1.313813658611069e+17, 1.31381365867982e+17, 1.31381365870482e+17, 1.313813658818883e+17, 1.313813658845445e+17, 1.313813658934508e+17, 1.313813658965757e+17, 1.313813659037632e+17, 1.313813659115757e+17, 1.313813659172008e+17, 1.313813659256381e+17, 1.313813659301695e+17, 1.313813659368882e+17, 1.313813659437632e+17, 1.313813659509508e+17, 1.31381365959232e+17, 1.313813659631383e+17, 1.313813659700132e+17, 1.313813659779821e+17, 1.313813659826694e+17, 1.313813659900132e+17, 1.313813659962633e+17, 1.313813660031383e+17, 1.31381366010482e+17, 1.313813660173569e+17, 1.313813660237632e+17, 1.313813660306382e+17, 1.313813660367319e+17, 1.31381366043607e+17, 1.31381366050482e+17, 1.313813660575132e+17, 1.313813660634508e+17, 1.313813660737632e+17, 1.31381366076107e+17, 1.313813660795444e+17, 1.313813660889196e+17, 1.313813660928259e+17, 1.31381366099857e+17, 1.313813661068883e+17, 1.31381366113607e+17, 1.313813661203258e+17, 1.313813661259507e+17, 1.313813661331383e+17, 1.31381366135482e+17, 1.313813661468883e+17, 1.313813661509508e+17, 1.313813661615758e+17, 1.313813661647008e+17, 1.31381366171732e+17, 1.313813661740756e+17, 1.313813661847008e+17, 1.31381366189857e+17, 1.313813661997007e+17, 1.313813662020444e+17, 1.31381366208607e+17, 1.313813662111069e+17, 1.313813662179821e+17, 1.313813662275132e+17, 1.313813662297007e+17, 1.313813662362633e+17, 1.31381366238607e+17, 1.313813662409507e+17, 1.313813662479821e+17, 1.313813662557946e+17, 1.313813662625133e+17, 1.313813662687633e+17, 1.313813662745445e+17, 1.313813662814195e+17, 1.313813662839195e+17, 1.31381366295482e+17, 1.313813662978257e+17, 1.313813663064195e+17, 1.313813663120444e+17, 1.313813663200133e+17, 1.313813663225133e+17, 1.313813663290757e+17, 1.313813663347008e+17, 1.313813663406382e+17, 1.313813663475132e+17, 1.313813663547008e+17, 1.31381366361732e+17, 1.313813663640758e+17, 1.313813663756383e+17, 1.31381366377982e+17, 1.313813663881382e+17, 1.31381366390482e+17, 1.313813663965757e+17, 1.313813664014195e+17, 1.313813664075133e+17, 1.313813664143882e+17, 1.31381366426732e+17, 1.313813664293883e+17, 1.313813664368883e+17, 1.31381366442982e+17, 1.313813664500133e+17, 1.313813664564195e+17, 1.313813664632945e+17, 1.313813664718883e+17, 1.31381366476107e+17, 1.313813664820444e+17, 1.313813664928257e+17, 1.313813664951695e+17, 1.313813665031383e+17, 1.31381366505482e+17, 1.313813665140758e+17, 1.313813665197007e+17, 1.313813665220445e+17, 1.313813665336069e+17, 1.313813665365757e+17, 1.313813665464195e+17, 1.313813665501695e+17, 1.313813665601695e+17, 1.313813665625133e+17, 1.31381366572357e+17, 1.313813665747008e+17, 1.313813665853257e+17, 1.313813665912632e+17, 1.313813665990757e+17, 1.313813666062633e+17, 1.313813666132945e+17, 1.313813666156383e+17, 1.313813666226696e+17, 1.313813666301695e+17, 1.31381366640482e+17, 1.313813666443882e+17, 1.313813666503256e+17, 1.313813666609508e+17, 1.313813666632945e+17, 1.313813666693883e+17, 1.313813666743882e+17, 1.313813666803258e+17, 1.313813666826696e+17, 1.313813666947007e+17, 1.313813667031383e+17, 1.313813667070446e+17, 1.313813667145445e+17, 1.313813667217321e+17, 1.313813667306382e+17, 1.31381366734857e+17, 1.313813667409508e+17, 1.313813667478258e+17, 1.31381366756732e+17, 1.313813667612632e+17, 1.313813667672008e+17, 1.313813667742319e+17, 1.313813667801695e+17, 1.31381366786732e+17, 1.313813667937632e+17, 1.313813668009507e+17, 1.313813668076695e+17, 1.313813668139195e+17, 1.313813668162632e+17, 1.313813668282945e+17, 1.313813668306382e+17, 1.313813668382945e+17, 1.313813668406383e+17, 1.313813668473571e+17, 1.313813668550132e+17, 1.31381366859232e+17, 1.313813668668883e+17, 1.31381366872357e+17, 1.313813668812632e+17, 1.313813668843882e+17, 1.31381366890482e+17, 1.31381366895482e+17, 1.313813668978258e+17, 1.313813669093883e+17, 1.313813669132945e+17, 1.313813669200132e+17, 1.313813669257946e+17, 1.31381366929857e+17, 1.313813669397007e+17, 1.313813669475132e+17, 1.313813669547007e+17, 1.31381366961732e+17, 1.313813669743884e+17, 1.313813669770445e+17, 1.313813669840758e+17, 1.31381366992982e+17, 1.313813669972008e+17, 1.313813670032945e+17, 1.313813670103258e+17, 1.313813670126696e+17, 1.313813670264195e+17, 1.31381367030482e+17, 1.313813670373569e+17, 1.313813670443882e+17, 1.31381367051732e+17, 1.313813670611069e+17, 1.313813670648571e+17, 1.313813670709508e+17, 1.31381367077982e+17, 1.313813670859507e+17, 1.313813670947008e+17, 1.31381367099232e+17, 1.313813671050132e+17, 1.313813671132945e+17, 1.313813671182945e+17, 1.313813671206382e+17, 1.313813671323571e+17, 1.313813671351695e+17, 1.313813671432945e+17, 1.313813671509508e+17, 1.313813671543882e+17, 1.313813671614195e+17, 1.313813671656383e+17, 1.313813671732945e+17, 1.313813671757944e+17, 1.313813671825133e+17, 1.31381367192357e+17, 1.313813671993883e+17, 1.313813672073571e+17, 1.313813672125133e+17, 1.313813672203258e+17, 1.313813672251695e+17, 1.313813672275132e+17, 1.313813672342319e+17, 1.31381367242357e+17, 1.313813672489196e+17, 1.313813672559507e+17, 1.313813672631383e+17, 1.313813672701696e+17, 1.313813672756383e+17, 1.313813672831383e+17, 1.313813672901695e+17, 1.313813672972008e+17, 1.313813673042321e+17, 1.313813673111071e+17, 1.31381367319232e+17, 1.313813673264195e+17, 1.313813673334508e+17, 1.313813673357946e+17, 1.313813673434508e+17, 1.313813673506382e+17, 1.313813673572008e+17, 1.313813673656383e+17, 1.313813673703258e+17, 1.313813673762632e+17, 1.313813673872008e+17, 1.31381367390482e+17, 1.313813673975132e+17, 1.313813674047008e+17, 1.313813674117321e+17, 1.313813674178258e+17, 1.313813674247008e+17, 1.313813674314195e+17, 1.313813674420445e+17, 1.313813674478257e+17, 1.313813674548571e+17, 1.313813674620444e+17, 1.313813674682945e+17, 1.313813674753257e+17, 1.313813674820444e+17, 1.313813674889196e+17, 1.313813674950132e+17, 1.313813675015758e+17, 1.313813675082945e+17, 1.313813675153257e+17, 1.313813675225133e+17, 1.313813675295446e+17, 1.313813675423571e+17, 1.313813675448571e+17, 1.313813675545445e+17, 1.313813675578257e+17, 1.313813675618883e+17, 1.31381367571732e+17, 1.313813675742319e+17, 1.313813675859507e+17, 1.313813675884508e+17, 1.313813675964196e+17, 1.313813676034508e+17, 1.313813676103258e+17, 1.31381367618607e+17, 1.313813676256383e+17, 1.31381367632357e+17, 1.313813676382945e+17, 1.31381367645482e+17, 1.313813676573571e+17, 1.313813676606382e+17, 1.313813676709508e+17, 1.313813676732945e+17, 1.313813676757944e+17, 1.313813676859507e+17, 1.313813676901695e+17, 1.313813676978258e+17, 1.313813677072008e+17, 1.31381367712357e+17, 1.313813677203258e+17, 1.313813677276695e+17, 1.313813677347008e+17, 1.313813677420444e+17, 1.313813677490757e+17, 1.313813677590757e+17, 1.313813677643882e+17, 1.313813677715757e+17, 1.31381367777982e+17, 1.313813677873571e+17, 1.31381367791732e+17, 1.313813677987633e+17, 1.313813678011071e+17, 1.313813678132945e+17, 1.313813678193883e+17, 1.31381367826107e+17, 1.313813678332945e+17, 1.313813678395446e+17, 1.313813678453257e+17, 1.313813678526694e+17, 1.313813678578258e+17, 1.313813678601695e+17, 1.313813678720444e+17, 1.31381367874857e+17, 1.31381367883607e+17, 1.313813678886071e+17, 1.313813678909508e+17, 1.313813679026696e+17, 1.31381367910482e+17, 1.313813679206382e+17, 1.313813679257946e+17, 1.313813679331383e+17, 1.313813679401695e+17, 1.313813679472008e+17, 1.313813679573571e+17, 1.31381367962357e+17, 1.313813679701695e+17, 1.313813679775132e+17, 1.313813679803258e+17, 1.313813679925133e+17, 1.313813680037632e+17, 1.31381368006107e+17, 1.313813680134508e+17, 1.313813680197007e+17, 1.31381368024857e+17, 1.313813680314195e+17, 1.31381368038607e+17, 1.313813680478258e+17, 1.313813680520445e+17, 1.31381368057982e+17, 1.313813680651695e+17, 1.313813680707945e+17, 1.313813680784507e+17, 1.313813680865757e+17, 1.313813680939195e+17, 1.313813680962632e+17, 1.313813681093883e+17, 1.31381368112982e+17, 1.313813681220445e+17, 1.313813681262633e+17, 1.313813681334508e+17, 1.313813681395446e+17, 1.313813681478257e+17, 1.313813681548571e+17, 1.313813681618883e+17, 1.313813681723571e+17, 1.31381368175482e+17, 1.313813681839195e+17, 1.313813681862633e+17, 1.313813681945444e+17, 1.313813681997007e+17, 1.313813682076695e+17, 1.313813682147007e+17, 1.313813682218883e+17, 1.313813682297007e+17, 1.313813682362633e+17, 1.313813682431382e+17, 1.313813682489196e+17, 1.31381368256107e+17, 1.313813682642321e+17, 1.313813682745445e+17, 1.313813682778257e+17, 1.313813682850132e+17, 1.313813682911069e+17, 1.313813682997007e+17, 1.313813683045444e+17, 1.313813683068882e+17, 1.313813683137632e+17, 1.313813683197007e+17, 1.313813683262633e+17, 1.31381368333607e+17, 1.313813683393883e+17, 1.313813683465757e+17, 1.313813683528257e+17, 1.313813683598569e+17, 1.313813683670445e+17, 1.313813683740758e+17, 1.313813683822007e+17, 1.313813683890757e+17, 1.313813683964195e+17, 1.31381368402357e+17, 1.313813684128257e+17, 1.313813684190757e+17, 1.313813684251695e+17, 1.313813684323571e+17, 1.313813684381382e+17, 1.313813684450132e+17, 1.313813684511069e+17, 1.313813684575132e+17, 1.313813684647008e+17, 1.31381368471732e+17, 1.313813684784508e+17, 1.313813684857946e+17, 1.313813684922007e+17, 1.313813685045445e+17, 1.313813685072008e+17, 1.313813685145445e+17, 1.313813685203258e+17, 1.313813685264195e+17, 1.313813685353257e+17, 1.313813685414195e+17, 1.31381368548607e+17, 1.313813685556383e+17, 1.313813685618883e+17, 1.313813685690757e+17, 1.313813685750132e+17, 1.313813685820444e+17, 1.313813685893883e+17, 1.313813685964196e+17, 1.31381368603607e+17, 1.313813686106382e+17, 1.313813686187633e+17, 1.31381368625482e+17, 1.313813686322008e+17, 1.313813686382945e+17, 1.313813686456383e+17, 1.313813686528257e+17, 1.313813686639195e+17, 1.313813686682945e+17, 1.313813686743882e+17, 1.313813686820445e+17, 1.313813686893883e+17, 1.31381368699857e+17, 1.313813687020445e+17, 1.313813687101695e+17, 1.313813687125133e+17, 1.313813687148571e+17, 1.313813687245445e+17, 1.313813687295446e+17, 1.31381368742357e+17, 1.313813687450132e+17, 1.313813687511069e+17, 1.313813687582945e+17, 1.313813687664195e+17, 1.313813687747008e+17, 1.313813687812632e+17, 1.31381368788607e+17, 1.313813687995444e+17, 1.313813688084508e+17, 1.313813688107945e+17, 1.313813688211071e+17, 1.313813688275132e+17, 1.313813688306382e+17, 1.313813688373569e+17, 1.313813688434508e+17, 1.313813688457944e+17, 1.313813688576695e+17, 1.313813688601695e+17, 1.313813688684507e+17, 1.313813688750132e+17, 1.313813688840758e+17, 1.313813688903258e+17, 1.313813688978258e+17, 1.313813689047007e+17, 1.313813689115757e+17, 1.313813689181382e+17, 1.313813689240758e+17, 1.313813689312632e+17, 1.31381368938607e+17, 1.313813689459507e+17, 1.313813689539195e+17, 1.313813689575132e+17, 1.313813689650132e+17, 1.31381368972357e+17, 1.313813689856383e+17, 1.31381368988607e+17, 1.313813689979821e+17, 1.31381369000482e+17, 1.31381369006107e+17, 1.313813690089196e+17, 1.31381369016107e+17, 1.31381369018607e+17, 1.313813690251695e+17, 1.313813690306382e+17, 1.313813690381382e+17, 1.313813690442321e+17, 1.313813690514195e+17, 1.313813690587633e+17, 1.31381369064857e+17, 1.313813690672008e+17, 1.31381369079232e+17, 1.313813690815757e+17, 1.313813690906382e+17, 1.313813690970445e+17, 1.313813691039195e+17, 1.313813691134508e+17, 1.313813691189196e+17, 1.31381369126107e+17, 1.313813691284507e+17, 1.313813691404819e+17, 1.31381369142982e+17, 1.313813691509508e+17, 1.313813691597007e+17, 1.313813691642319e+17, 1.313813691703258e+17, 1.313813691776695e+17, 1.31381369184857e+17, 1.313813691918883e+17, 1.313813691987633e+17, 1.313813692076695e+17, 1.31381369211732e+17, 1.313813692173571e+17, 1.31381369225482e+17, 1.313813692315757e+17, 1.313813692339195e+17, 1.313813692447008e+17, 1.313813692484508e+17, 1.31381369255482e+17, 1.313813692628257e+17, 1.31381369271732e+17, 1.313813692762633e+17, 1.313813692839195e+17, 1.313813692931383e+17, 1.313813692965757e+17, 1.313813693026694e+17, 1.31381369309857e+17, 1.31381369316732e+17, 1.313813693234508e+17, 1.313813693295444e+17, 1.31381369336107e+17, 1.313813693434508e+17, 1.313813693506382e+17, 1.313813693573569e+17, 1.313813693672008e+17, 1.313813693711069e+17, 1.31381369377982e+17, 1.313813693804819e+17, 1.313813693914194e+17, 1.31381369397982e+17, 1.313813694051695e+17, 1.313813694140758e+17, 1.313813694189196e+17, 1.313813694250132e+17, 1.313813694309507e+17, 1.313813694378258e+17, 1.313813694401695e+17, 1.313813694518883e+17, 1.313813694543882e+17, 1.313813694650132e+17, 1.313813694722007e+17, 1.313813694776695e+17, 1.313813694839195e+17, 1.313813694911069e+17, 1.313813694993883e+17, 1.313813695059507e+17, 1.31381369513607e+17, 1.31381369520482e+17, 1.313813695275132e+17, 1.313813695347007e+17, 1.313813695420444e+17, 1.313813695539195e+17, 1.313813695573569e+17, 1.313813695642321e+17, 1.313813695706382e+17, 1.313813695775133e+17, 1.313813695848571e+17, 1.313813695922007e+17, 1.313813695995444e+17, 1.313813696054821e+17, 1.313813696128257e+17, 1.313813696201696e+17, 1.313813696272008e+17, 1.313813696342321e+17, 1.313813696418883e+17, 1.313813696515758e+17, 1.313813696540758e+17, 1.31381369661732e+17, 1.313813696681382e+17, 1.313813696762632e+17, 1.313813696836069e+17, 1.313813696915757e+17, 1.31381369698607e+17, 1.313813697057946e+17, 1.31381369712982e+17, 1.31381369719232e+17, 1.313813697257946e+17, 1.313813697348571e+17, 1.313813697397009e+17, 1.313813697467319e+17, 1.313813697537633e+17, 1.313813697612632e+17, 1.31381369768607e+17, 1.313813697753257e+17, 1.313813697826694e+17, 1.313813697889196e+17, 1.313813697981382e+17, 1.313813698032945e+17, 1.313813698104819e+17, 1.313813698182945e+17, 1.313813698240758e+17, 1.313813698264195e+17, 1.313813698387633e+17, 1.313813698415757e+17, 1.313813698512632e+17, 1.313813698550132e+17, 1.313813698620445e+17, 1.313813698703258e+17, 1.313813698762632e+17, 1.313813698850132e+17, 1.313813698890757e+17, 1.313813698914195e+17, 1.313813699037633e+17, 1.313813699089196e+17, 1.31381369915482e+17, 1.313813699222007e+17, 1.313813699348571e+17, 1.313813699372008e+17, 1.313813699432946e+17, 1.313813699476695e+17, 1.31381369953607e+17, 1.313813699607945e+17, 1.313813699725133e+17, 1.313813699748571e+17, 1.313813699772008e+17, 1.31381369986107e+17, 1.313813699904819e+17, 1.313813699973571e+17, 1.313813700045445e+17, 1.31381370013607e+17, 1.313813700172008e+17, 1.313813700264196e+17, 1.313813700304819e+17, 1.313813700372006e+17, 1.313813700445445e+17, 1.31381370052982e+17, 1.313813700611071e+17, 1.313813700682945e+17, 1.313813700751695e+17, 1.313813700809508e+17, 1.31381370087982e+17, 1.313813700950132e+17, 1.31381370102357e+17, 1.31381370112357e+17, 1.313813701176695e+17, 1.313813701248571e+17, 1.313813701301695e+17, 1.313813701368882e+17, 1.313813701443882e+17, 1.31381370151732e+17, 1.313813701578258e+17, 1.313813701647007e+17, 1.313813701717321e+17, 1.313813701789196e+17, 1.31381370186107e+17, 1.313813701932945e+17, 1.313813702014195e+17, 1.313813702072008e+17, 1.313813702153258e+17, 1.313813702176695e+17, 1.313813702275133e+17, 1.313813702325133e+17, 1.313813702407945e+17, 1.313813702481382e+17, 1.313813702511069e+17, 1.313813702631383e+17, 1.313813702714195e+17, 1.313813702768883e+17, 1.313813702839195e+17, 1.313813702911069e+17, 1.313813702973571e+17, 1.313813703045445e+17, 1.313813703114195e+17, 1.313813703175132e+17, 1.313813703257944e+17, 1.313813703378257e+17, 1.313813703411071e+17, 1.313813703470445e+17, 1.313813703540758e+17, 1.31381370362357e+17, 1.31381370369857e+17, 1.313813703787633e+17, 1.313813703822007e+17, 1.313813703889194e+17, 1.313813703943882e+17, 1.31381370396732e+17, 1.313813704090757e+17, 1.313813704139195e+17, 1.313813704162632e+17, 1.313813704222007e+17, 1.313813704322007e+17, 1.313813704345445e+17, 1.313813704472008e+17, 1.31381370453607e+17, 1.313813704637632e+17, 1.313813704668883e+17, 1.313813704748571e+17, 1.31381370478607e+17, 1.31381370484857e+17, 1.313813704918883e+17, 1.31381370499232e+17, 1.31381370506107e+17, 1.313813705128257e+17, 1.313813705200132e+17, 1.31381370526732e+17, 1.313813705334508e+17, 1.313813705403258e+17, 1.313813705478258e+17, 1.313813705547008e+17, 1.313813705622007e+17, 1.313813705700132e+17, 1.31381370577982e+17, 1.313813705823571e+17, 1.313813705897009e+17, 1.313813705967319e+17, 1.313813706031383e+17, 1.313813706103258e+17, 1.313813706176695e+17, 1.313813706247007e+17, 1.313813706318883e+17, 1.313813706393883e+17, 1.313813706420445e+17, 1.313813706545445e+17, 1.313813706606383e+17, 1.313813706686071e+17, 1.31381370675482e+17, 1.313813706790757e+17, 1.31381370686732e+17, 1.313813706943882e+17, 1.313813707015757e+17, 1.313813707095444e+17, 1.313813707145444e+17, 1.313813707170445e+17, 1.313813707287633e+17, 1.313813707339195e+17, 1.313813707412632e+17, 1.313813707484507e+17, 1.313813707554821e+17, 1.313813707626694e+17, 1.313813707695446e+17, 1.313813707776695e+17, 1.313813707847008e+17, 1.313813707918883e+17, 1.313813707989196e+17, 1.313813708056383e+17, 1.313813708118883e+17, 1.313813708187633e+17, 1.31381370825482e+17, 1.31381370832357e+17, 1.313813708414195e+17, 1.31381370846107e+17, 1.31381370855482e+17, 1.313813708606382e+17, 1.313813708648571e+17, 1.31381370874857e+17, 1.313813708828257e+17, 1.313813708900132e+17, 1.313813708972008e+17, 1.313813709051695e+17, 1.313813709073571e+17, 1.31381370919232e+17, 1.313813709215757e+17, 1.313813709332945e+17, 1.313813709356383e+17, 1.313813709462633e+17, 1.313813709495444e+17, 1.31381370956107e+17, 1.313813709620445e+17, 1.313813709720444e+17, 1.313813709759508e+17, 1.313813709839196e+17, 1.313813709889196e+17, 1.313813710022008e+17, 1.313813710043882e+17, 1.313813710103258e+17, 1.313813710153257e+17, 1.313813710231382e+17, 1.313813710312634e+17, 1.313813710386071e+17, 1.313813710432945e+17, 1.313813710507945e+17, 1.313813710579821e+17, 1.313813710651695e+17, 1.31381371072357e+17, 1.313813710747008e+17, 1.313813710868882e+17, 1.313813710942319e+17, 1.313813710989196e+17, 1.313813711031383e+17, 1.313813711131382e+17, 1.31381371115482e+17, 1.313813711276695e+17, 1.313813711347008e+17, 1.313813711420444e+17, 1.313813711475132e+17, 1.313813711545445e+17, 1.31381371163607e+17, 1.31381371169857e+17, 1.313813711770445e+17, 1.313813711834508e+17, 1.313813711897007e+17, 1.313813711964195e+17, 1.313813712025133e+17, 1.313813712100133e+17, 1.313813712182945e+17, 1.313813712237632e+17, 1.31381371226107e+17, 1.313813712390757e+17, 1.313813712439196e+17, 1.313813712525133e+17, 1.313813712606382e+17, 1.313813712681382e+17, 1.313813712751695e+17, 1.313813712775132e+17, 1.313813712893883e+17, 1.313813712950132e+17, 1.313813713012632e+17, 1.31381371303607e+17, 1.313813713157944e+17, 1.313813713211071e+17, 1.313813713272008e+17, 1.313813713342319e+17, 1.313813713414195e+17, 1.31381371348607e+17, 1.31381371354857e+17, 1.313813713617321e+17, 1.313813713640758e+17, 1.313813713759507e+17, 1.313813713782945e+17, 1.313813713862633e+17, 1.313813713934508e+17, 1.313813714004819e+17, 1.313813714072008e+17, 1.313813714142321e+17, 1.313813714203258e+17, 1.313813714272008e+17, 1.313813714342319e+17, 1.313813714409508e+17, 1.313813714497007e+17, 1.313813714550132e+17, 1.31381371462357e+17, 1.313813714695444e+17, 1.313813714765757e+17, 1.313813714859507e+17, 1.313813714907945e+17, 1.31381371497982e+17, 1.31381371504857e+17, 1.313813715107945e+17, 1.313813715178258e+17, 1.31381371529857e+17, 1.31381371532982e+17, 1.313813715400133e+17, 1.31381371542357e+17, 1.313813715484508e+17, 1.313813715557944e+17, 1.313813715647008e+17, 1.313813715706382e+17, 1.313813715778257e+17, 1.313813715840758e+17, 1.313813715914195e+17, 1.313813715984507e+17, 1.313813716065757e+17, 1.313813716118883e+17, 1.313813716170445e+17, 1.31381371626732e+17, 1.313813716340758e+17, 1.31381371642357e+17, 1.313813716500133e+17, 1.313813716562632e+17, 1.313813716645445e+17, 1.31381371677982e+17, 1.313813716803258e+17, 1.313813716864195e+17, 1.313813716922008e+17, 1.31381371699857e+17, 1.31381371709232e+17, 1.313813717125133e+17, 1.31381371718607e+17, 1.313813717293883e+17, 1.313813717326694e+17, 1.31381371739857e+17, 1.313813717462633e+17, 1.313813717531383e+17, 1.313813717595444e+17, 1.313813717656383e+17, 1.313813717747007e+17, 1.313813717822008e+17, 1.313813717889196e+17, 1.313813717959507e+17, 1.313813718037632e+17, 1.313813718114195e+17, 1.313813718211071e+17, 1.313813718248571e+17, 1.313813718312632e+17, 1.313813718382945e+17, 1.313813718470445e+17, 1.31381371851732e+17, 1.313813718540758e+17, 1.313813718657944e+17, 1.31381371869232e+17, 1.313813718787633e+17, 1.313813718822007e+17, 1.313813718847007e+17, 1.313813718953257e+17, 1.313813719034508e+17, 1.313813719107945e+17, 1.313813719168882e+17, 1.31381371919232e+17, 1.313813719248571e+17, 1.313813719326694e+17, 1.31381371939232e+17, 1.31381371946107e+17, 1.313813719545445e+17, 1.313813719597007e+17, 1.313813719665757e+17, 1.313813719739195e+17, 1.313813719811069e+17, 1.313813719884507e+17, 1.31381371995482e+17, 1.313813720025133e+17, 1.313813720093883e+17, 1.313813720154821e+17, 1.313813720214195e+17, 1.313813720293883e+17, 1.313813720340756e+17, 1.313813720420444e+17, 1.313813720470445e+17, 1.31381372055482e+17, 1.313813720626694e+17, 1.313813720695446e+17, 1.313813720776695e+17, 1.313813720839195e+17, 1.313813720887633e+17, 1.31381372095482e+17, 1.313813721023571e+17, 1.313813721132945e+17, 1.313813721159507e+17, 1.313813721225133e+17, 1.313813721278258e+17, 1.313813721340758e+17, 1.313813721409507e+17, 1.313813721432945e+17, 1.313813721550132e+17, 1.313813721575132e+17, 1.313813721682945e+17, 1.31381372172357e+17, 1.313813721820445e+17, 1.313813721872006e+17, 1.313813721943882e+17, 1.313813722011069e+17, 1.313813722079821e+17, 1.313813722137632e+17, 1.313813722214195e+17, 1.313813722314195e+17, 1.313813722376695e+17, 1.313813722412632e+17, 1.313813722481382e+17, 1.313813722550132e+17, 1.313813722620445e+17, 1.313813722684507e+17, 1.313813722757944e+17, 1.31381372284857e+17, 1.313813722928257e+17, 1.31381372295482e+17, 1.313813723025133e+17, 1.313813723072008e+17, 1.313813723153257e+17, 1.313813723200133e+17, 1.313813723262633e+17, 1.313813723340758e+17, 1.313813723387633e+17, 1.31381372346107e+17, 1.313813723534508e+17, 1.313813723595444e+17, 1.313813723668882e+17, 1.313813723768883e+17, 1.313813723822007e+17, 1.31381372389232e+17, 1.313813723915758e+17, 1.31381372403607e+17, 1.313813724059507e+17, 1.313813724172008e+17, 1.313813724195444e+17, 1.313813724218883e+17, 1.313813724315758e+17, 1.313813724357946e+17, 1.31381372442982e+17, 1.313813724537632e+17, 1.313813724562632e+17, 1.313813724625133e+17, 1.313813724686071e+17, 1.31381372476107e+17, 1.313813724832945e+17, 1.313813724856383e+17, 1.313813724964195e+17, 1.31381372502982e+17, 1.31381372509232e+17, 1.313813725164195e+17, 1.313813725215757e+17, 1.313813725301695e+17, 1.313813725325133e+17, 1.313813725395444e+17, 1.313813725451695e+17, 1.313813725532945e+17, 1.313813725587633e+17, 1.313813725611071e+17, 1.313813725732945e+17, 1.313813725789196e+17, 1.313813725812632e+17, 1.313813725932945e+17, 1.313813725956383e+17, 1.313813726057944e+17, 1.313813726103258e+17, 1.313813726193883e+17, 1.313813726231383e+17, 1.313813726300132e+17, 1.31381372635482e+17, 1.313813726426696e+17, 1.313813726500132e+17, 1.313813726526696e+17, 1.313813726653257e+17, 1.313813726707945e+17, 1.31381372679232e+17, 1.313813726864195e+17, 1.313813726934508e+17, 1.313813726998569e+17, 1.313813727068883e+17, 1.313813727150132e+17, 1.31381372722357e+17, 1.313813727293883e+17, 1.31381372739232e+17, 1.313813727431383e+17, 1.313813727495444e+17, 1.31381372756732e+17, 1.313813727632946e+17, 1.313813727714195e+17, 1.313813727797009e+17, 1.313813727867319e+17, 1.313813727932945e+17, 1.313813727993883e+17, 1.313813728064196e+17, 1.313813728137633e+17, 1.313813728206382e+17, 1.313813728289196e+17, 1.313813728359507e+17, 1.31381372842982e+17, 1.313813728509508e+17, 1.31381372856107e+17, 1.313813728648571e+17, 1.313813728695446e+17, 1.313813728764195e+17, 1.31381372883607e+17, 1.31381372889857e+17, 1.313813728990757e+17, 1.313813729043882e+17, 1.313813729115758e+17, 1.313813729218883e+17, 1.313813729242321e+17, 1.313813729314195e+17, 1.313813729362632e+17, 1.313813729434508e+17, 1.313813729506382e+17, 1.313813729576695e+17, 1.313813729622007e+17, 1.313813729692321e+17, 1.313813729756383e+17, 1.313813729801695e+17, 1.313813729872008e+17, 1.313813729945445e+17, 1.31381373001732e+17, 1.313813730100133e+17, 1.313813730154821e+17, 1.313813730215758e+17, 1.31381373028607e+17, 1.313813730364195e+17, 1.313813730415758e+17, 1.313813730489196e+17, 1.31381373056107e+17, 1.313813730645445e+17, 1.313813730707945e+17, 1.313813730731383e+17, 1.31381373086107e+17, 1.313813730931383e+17, 1.313813730997007e+17, 1.313813731018883e+17, 1.313813731139195e+17, 1.313813731212632e+17, 1.313813731284508e+17, 1.313813731359507e+17, 1.313813731420444e+17, 1.313813731503258e+17, 1.313813731576695e+17, 1.313813731645444e+17, 1.313813731668882e+17, 1.313813731789196e+17, 1.313813731812634e+17, 1.31381373190482e+17, 1.313813731965757e+17, 1.313813732034508e+17, 1.313813732084507e+17, 1.31381373215482e+17, 1.313813732222007e+17, 1.313813732309508e+17, 1.313813732370445e+17, 1.313813732440756e+17, 1.313813732514195e+17, 1.313813732614195e+17, 1.313813732664196e+17, 1.313813732734508e+17, 1.313813732868883e+17, 1.313813732893883e+17, 1.313813732950132e+17, 1.313813732978258e+17, 1.313813733043882e+17, 1.313813733106383e+17, 1.313813733178258e+17, 1.313813733206382e+17, 1.313813733301696e+17, 1.313813733376695e+17, 1.313813733437632e+17, 1.313813733507945e+17, 1.31381373356732e+17, 1.313813733637632e+17, 1.31381373376732e+17, 1.313813733790757e+17, 1.313813733814195e+17, 1.313813733903258e+17, 1.31381373394857e+17, 1.313813734050132e+17, 1.313813734076695e+17, 1.313813734156383e+17, 1.313813734203258e+17, 1.313813734306382e+17, 1.31381373432982e+17, 1.313813734420444e+17, 1.313813734451695e+17, 1.313813734475132e+17, 1.31381373459232e+17, 1.313813734643884e+17, 1.31381373466732e+17, 1.313813734734509e+17, 1.313813734797007e+17, 1.313813734856383e+17, 1.313813734931383e+17, 1.313813735003258e+17, 1.313813735076695e+17, 1.313813735176695e+17, 1.313813735256383e+17, 1.313813735312632e+17, 1.313813735364195e+17, 1.313813735447008e+17, 1.313813735522007e+17, 1.313813735595444e+17, 1.313813735665757e+17, 1.313813735731383e+17, 1.313813735765757e+17, 1.31381373586107e+17, 1.313813735940758e+17, 1.313813736022008e+17, 1.313813736093882e+17, 1.31381373616732e+17, 1.313813736239195e+17, 1.313813736314195e+17, 1.313813736393883e+17, 1.313813736465757e+17, 1.313813736495444e+17, 1.313813736617321e+17, 1.313813736682944e+17, 1.313813736751695e+17, 1.313813736826696e+17, 1.313813736900133e+17, 1.31381373696107e+17, 1.313813737045445e+17, 1.313813737128257e+17, 1.313813737200133e+17, 1.313813737273571e+17, 1.31381373733607e+17, 1.313813737414195e+17, 1.313813737489194e+17, 1.313813737559508e+17, 1.313813737584508e+17, 1.313813737712632e+17, 1.313813737775132e+17, 1.313813737837632e+17, 1.313813737901695e+17, 1.313813737978258e+17, 1.31381373803607e+17, 1.313813738106383e+17, 1.313813738178258e+17, 1.313813738232945e+17, 1.313813738306383e+17, 1.313813738378257e+17, 1.31381373845482e+17, 1.31381373855482e+17, 1.313813738579821e+17, 1.313813738651695e+17, 1.313813738718883e+17, 1.313813738812632e+17, 1.31381373886732e+17, 1.313813738939195e+17, 1.313813739012632e+17, 1.313813739082945e+17, 1.313813739173569e+17, 1.313813739231383e+17, 1.313813739334508e+17, 1.313813739378257e+17, 1.313813739456383e+17, 1.313813739542319e+17, 1.313813739593883e+17, 1.31381373961732e+17, 1.313813739743882e+17, 1.313813739797007e+17, 1.313813739856383e+17, 1.313813739931382e+17, 1.313813740028257e+17, 1.313813740065757e+17, 1.313813740142321e+17, 1.313813740222008e+17, 1.31381374027982e+17, 1.313813740350132e+17, 1.313813740375132e+17, 1.313813740445445e+17, 1.31381374052357e+17, 1.313813740600133e+17, 1.31381374064857e+17, 1.313813740720444e+17, 1.313813740775132e+17, 1.313813740850132e+17, 1.31381374092357e+17, 1.313813740964195e+17, 1.31381374105482e+17, 1.313813741126696e+17, 1.31381374119857e+17, 1.313813741273569e+17, 1.313813741336069e+17, 1.313813741417321e+17, 1.313813741476695e+17, 1.313813741557946e+17, 1.31381374162357e+17, 1.313813741697007e+17, 1.313813741768883e+17, 1.313813741847007e+17, 1.313813741886071e+17, 1.313813741970445e+17, 1.313813742032945e+17, 1.313813742081382e+17, 1.313813742140758e+17, 1.313813742218883e+17, 1.313813742318883e+17, 1.313813742345445e+17, 1.313813742368882e+17, 1.313813742490757e+17, 1.313813742525133e+17, 1.313813742604819e+17, 1.313813742701695e+17, 1.313813742762632e+17, 1.31381374284857e+17, 1.313813742922007e+17, 1.313813742990758e+17, 1.313813743109508e+17, 1.313813743143882e+17, 1.313813743228257e+17, 1.313813743281382e+17, 1.313813743356383e+17, 1.313813743420444e+17, 1.31381374345482e+17, 1.313813743573571e+17, 1.313813743643882e+17, 1.313813743726696e+17, 1.31381374379857e+17, 1.313813743862632e+17, 1.313813743907945e+17, 1.313813744007945e+17, 1.313813744107945e+17, 1.313813744143882e+17, 1.313813744167319e+17, 1.313813744293883e+17, 1.313813744334508e+17, 1.313813744406383e+17, 1.313813744479821e+17, 1.313813744542321e+17, 1.313813744628257e+17, 1.313813744711071e+17, 1.31381374478607e+17, 1.313813744857944e+17, 1.313813744881382e+17, 1.31381374500482e+17, 1.313813745050134e+17, 1.313813745131382e+17, 1.313813745203258e+17, 1.31381374526107e+17, 1.313813745337633e+17, 1.313813745401695e+17, 1.313813745476695e+17, 1.313813745542321e+17, 1.313813745615758e+17, 1.313813745678257e+17, 1.313813745753257e+17, 1.313813745822008e+17, 1.313813745862632e+17, 1.313813745957944e+17, 1.313813746031383e+17, 1.313813746125133e+17, 1.313813746201695e+17, 1.31381374626732e+17, 1.31381374632982e+17, 1.31381374640482e+17, 1.31381374648607e+17, 1.313813746556383e+17, 1.31381374662982e+17, 1.31381374672982e+17, 1.313813746765757e+17, 1.31381374683607e+17, 1.313813746906382e+17, 1.31381374699232e+17, 1.313813747059507e+17, 1.313813747176695e+17, 1.313813747209508e+17, 1.313813747268882e+17, 1.313813747347008e+17, 1.313813747432945e+17, 1.31381374751732e+17, 1.313813747582945e+17, 1.313813747611069e+17, 1.31381374773607e+17, 1.313813747803258e+17, 1.313813747876695e+17, 1.313813747950132e+17, 1.31381374802357e+17, 1.313813748095444e+17, 1.313813748170445e+17, 1.31381374822357e+17, 1.313813748325133e+17, 1.31381374842357e+17, 1.313813748462632e+17, 1.313813748534508e+17, 1.313813748618883e+17, 1.313813748728257e+17, 1.31381374875482e+17, 1.313813748826694e+17, 1.313813748887631e+17, 1.313813748970445e+17, 1.313813749042321e+17, 1.313813749122008e+17, 1.313813749193883e+17, 1.313813749314195e+17, 1.31381374934857e+17, 1.313813749428257e+17, 1.313813749484508e+17, 1.313813749575132e+17, 1.313813749615757e+17, 1.313813749639195e+17, 1.313813749762632e+17, 1.313813749790757e+17, 1.31381374986107e+17, 1.313813749925133e+17, 1.313813750015757e+17, 1.313813750062633e+17, 1.313813750139195e+17, 1.313813750215758e+17, 1.313813750290757e+17, 1.313813750365757e+17, 1.31381375044857e+17, 1.313813750512632e+17, 1.313813750587633e+17, 1.313813750662633e+17, 1.313813750734508e+17, 1.313813750856383e+17, 1.31381375089232e+17, 1.313813750976695e+17, 1.313813751022008e+17, 1.313813751147008e+17, 1.313813751181382e+17, 1.31381375123607e+17, 1.313813751322007e+17, 1.313813751411071e+17, 1.313813751447008e+17, 1.313813751522007e+17, 1.313813751575133e+17, 1.313813751648571e+17, 1.313813751736069e+17, 1.313813751818883e+17, 1.313813751893882e+17, 1.313813751973569e+17, 1.313813751997007e+17, 1.313813752109508e+17, 1.313813752181382e+17, 1.313813752253257e+17, 1.313813752328257e+17, 1.31381375239232e+17, 1.313813752475132e+17, 1.31381375255482e+17, 1.313813752653257e+17, 1.313813752700133e+17, 1.31381375276732e+17, 1.313813752839195e+17, 1.313813752922007e+17, 1.313813753020445e+17, 1.31381375306107e+17, 1.313813753147008e+17, 1.31381375319857e+17, 1.313813753222008e+17, 1.313813753347007e+17, 1.313813753403258e+17, 1.313813753462632e+17, 1.313813753554821e+17, 1.313813753626694e+17, 1.31381375369232e+17, 1.313813753765756e+17, 1.313813753868882e+17, 1.31381375389232e+17, 1.313813753915758e+17, 1.313813754007945e+17, 1.31381375404857e+17, 1.313813754111069e+17, 1.313813754182945e+17, 1.313813754257944e+17, 1.313813754343882e+17, 1.313813754425133e+17, 1.313813754522007e+17, 1.313813754562633e+17, 1.31381375458607e+17, 1.313813754707945e+17, 1.313813754756383e+17, 1.313813754845445e+17, 1.313813754873571e+17, 1.31381375494857e+17, 1.313813754997007e+17, 1.31381375506107e+17, 1.31381375513607e+17, 1.313813755220445e+17, 1.313813755275133e+17, 1.313813755376695e+17, 1.313813755428257e+17, 1.31381375550482e+17, 1.313813755587633e+17, 1.313813755650132e+17, 1.313813755717321e+17, 1.31381375578607e+17, 1.313813755868883e+17, 1.313813755942321e+17, 1.313813755982944e+17, 1.313813756057946e+17, 1.313813756182945e+17, 1.313813756220444e+17, 1.313813756282945e+17, 1.313813756356383e+17, 1.31381375642357e+17, 1.313813756497007e+17, 1.313813756553257e+17, 1.313813756626694e+17, 1.313813756682945e+17, 1.313813756753257e+17, 1.313813756845444e+17, 1.313813756893883e+17, 1.313813756975133e+17, 1.313813757047007e+17, 1.313813757120445e+17, 1.31381375719857e+17, 1.31381375726107e+17, 1.313813757332945e+17, 1.313813757406383e+17, 1.313813757489194e+17, 1.313813757547008e+17, 1.313813757629819e+17, 1.313813757703258e+17, 1.313813757773571e+17, 1.31381375785482e+17, 1.313813757920444e+17, 1.313813757993883e+17, 1.31381375806732e+17, 1.313813758137632e+17, 1.313813758206382e+17, 1.313813758282945e+17, 1.313813758353257e+17, 1.31381375842357e+17, 1.313813758506383e+17, 1.313813758589194e+17, 1.313813758673569e+17, 1.313813758742321e+17, 1.313813758815758e+17, 1.313813758872008e+17, 1.313813758957946e+17, 1.313813759032945e+17, 1.313813759095446e+17, 1.313813759173571e+17, 1.313813759234508e+17, 1.313813759257944e+17, 1.313813759384507e+17, 1.313813759443882e+17, 1.31381375951732e+17, 1.313813759590757e+17, 1.313813759668883e+17, 1.313813759712632e+17, 1.313813759770445e+17, 1.313813759847007e+17, 1.313813759932945e+17, 1.313813759975132e+17, 1.313813760040758e+17, 1.313813760114195e+17, 1.313813760178258e+17, 1.313813760250132e+17, 1.313813760325133e+17, 1.313813760420445e+17, 1.313813760478257e+17, 1.313813760514195e+17, 1.313813760622008e+17, 1.313813760693883e+17, 1.313813760768883e+17, 1.313813760850132e+17, 1.313813760914195e+17, 1.31381376098607e+17, 1.31381376106107e+17, 1.313813761084508e+17, 1.313813761150132e+17, 1.313813761212632e+17, 1.313813761301695e+17, 1.31381376135482e+17, 1.313813761437632e+17, 1.313813761512632e+17, 1.313813761584507e+17, 1.313813761668882e+17, 1.313813761745445e+17, 1.313813761828257e+17, 1.313813761900132e+17, 1.313813761973569e+17, 1.313813762037633e+17, 1.313813762089194e+17, 1.313813762112632e+17, 1.313813762239195e+17, 1.31381376229232e+17, 1.313813762315758e+17, 1.313813762439195e+17, 1.313813762473571e+17, 1.313813762497007e+17, 1.313813762622007e+17, 1.313813762697007e+17, 1.313813762720444e+17, 1.313813762847007e+17, 1.313813762886071e+17, 1.31381376299857e+17, 1.313813763031383e+17, 1.313813763100133e+17, 1.313813763164195e+17, 1.313813763226696e+17, 1.31381376329857e+17, 1.313813763373571e+17, 1.313813763451695e+17, 1.31381376352357e+17, 1.313813763597007e+17, 1.313813763662632e+17, 1.31381376373607e+17, 1.313813763787633e+17, 1.313813763873569e+17, 1.313813763945445e+17, 1.313813764028259e+17, 1.313813764112632e+17, 1.313813764186071e+17, 1.31381376425482e+17, 1.31381376432982e+17, 1.313813764400133e+17, 1.313813764522007e+17, 1.313813764547008e+17, 1.313813764618883e+17, 1.313813764687633e+17, 1.313813764757946e+17, 1.313813764781382e+17, 1.313813764903258e+17, 1.31381376494857e+17, 1.31381376502357e+17, 1.313813765089196e+17, 1.313813765204819e+17, 1.31381376522982e+17, 1.313813765314195e+17, 1.313813765362632e+17, 1.313813765434508e+17, 1.313813765545445e+17, 1.313813765572008e+17, 1.313813765645445e+17, 1.313813765709508e+17, 1.313813765782945e+17, 1.313813765856383e+17, 1.313813765928257e+17, 1.313813766011069e+17, 1.313813766082945e+17, 1.313813766173571e+17, 1.313813766237632e+17, 1.31381376632982e+17, 1.313813766393883e+17, 1.313813766465757e+17, 1.313813766553257e+17, 1.31381376659232e+17, 1.313813766697007e+17, 1.313813766781382e+17, 1.313813766814195e+17, 1.313813766839195e+17, 1.313813766943882e+17, 1.313813766984507e+17, 1.313813767078258e+17, 1.313813767122007e+17, 1.313813767145445e+17, 1.313813767254821e+17, 1.313813767322008e+17, 1.313813767395446e+17, 1.31381376746732e+17, 1.313813767539195e+17, 1.313813767597007e+17, 1.313813767670445e+17, 1.313813767745445e+17, 1.313813767809508e+17, 1.313813767872006e+17, 1.313813767942321e+17, 1.313813768003258e+17, 1.313813768075132e+17, 1.313813768147008e+17, 1.313813768220445e+17, 1.313813768317321e+17, 1.313813768359508e+17, 1.313813768382945e+17, 1.313813768503256e+17, 1.313813768607945e+17, 1.313813768640758e+17, 1.313813768709508e+17, 1.313813768787633e+17, 1.313813768857946e+17, 1.31381376892982e+17, 1.313813769031383e+17, 1.313813769073569e+17, 1.313813769136069e+17, 1.313813769209508e+17, 1.313813769275132e+17, 1.313813769364196e+17, 1.313813769403258e+17, 1.313813769472008e+17, 1.313813769553257e+17, 1.313813769628257e+17, 1.313813769709508e+17, 1.313813769732945e+17, 1.313813769859507e+17, 1.313813769914195e+17, 1.313813769939195e+17, 1.313813770015757e+17, 1.313813770118883e+17, 1.313813770156381e+17, 1.313813770226696e+17, 1.313813770311071e+17, 1.313813770401696e+17, 1.313813770457946e+17, 1.31381377053607e+17, 1.31381377059857e+17, 1.313813770676695e+17, 1.313813770750132e+17, 1.313813770822007e+17, 1.313813770890757e+17, 1.31381377096732e+17, 1.313813771039196e+17, 1.313813771073569e+17, 1.313813771182944e+17, 1.313813771262632e+17, 1.31381377133607e+17, 1.313813771409508e+17, 1.313813771432945e+17, 1.313813771557944e+17, 1.313813771595444e+17, 1.313813771618883e+17, 1.313813771731383e+17, 1.313813771787633e+17, 1.313813771851694e+17, 1.313813771925133e+17, 1.313813772000133e+17, 1.313813772056383e+17, 1.313813772142319e+17, 1.313813772165757e+17, 1.31381377228607e+17, 1.313813772309508e+17, 1.313813772426696e+17, 1.313813772450132e+17, 1.313813772526696e+17, 1.313813772570445e+17, 1.313813772651695e+17, 1.313813772781382e+17, 1.31381377280482e+17, 1.31381377286107e+17, 1.313813772931382e+17, 1.313813773003258e+17, 1.313813773075133e+17, 1.313813773159508e+17, 1.313813773232945e+17, 1.313813773315757e+17, 1.313813773384508e+17, 1.313813773456383e+17, 1.313813773489196e+17, 1.313813773576695e+17, 1.313813773659507e+17, 1.313813773722007e+17, 1.313813773790758e+17, 1.31381377385482e+17, 1.313813773922007e+17, 1.313813773997007e+17, 1.31381377406107e+17, 1.313813774134508e+17, 1.313813774234508e+17, 1.313813774276695e+17, 1.313813774345445e+17, 1.313813774415757e+17, 1.313813774501696e+17, 1.313813774565757e+17, 1.313813774637633e+17, 1.313813774709508e+17, 1.313813774784507e+17, 1.31381377485482e+17, 1.313813774965757e+17, 1.313813775003258e+17, 1.313813775131382e+17, 1.313813775159507e+17, 1.31381377525482e+17, 1.313813775301695e+17, 1.313813775372008e+17, 1.313813775443884e+17, 1.313813775515758e+17, 1.313813775584508e+17, 1.313813775637633e+17, 1.313813775701695e+17, 1.31381377578607e+17, 1.31381377584857e+17, 1.31381377592982e+17, 1.313813775997009e+17, 1.313813776051695e+17, 1.313813776132945e+17, 1.313813776195444e+17, 1.313813776265757e+17, 1.31381377633607e+17, 1.313813776411069e+17, 1.313813776512632e+17, 1.313813776565757e+17, 1.313813776637632e+17, 1.31381377666107e+17, 1.313813776778257e+17, 1.31381377681732e+17, 1.313813776945445e+17, 1.313813776972008e+17, 1.313813777042321e+17, 1.313813777107945e+17, 1.313813777184507e+17, 1.31381377725482e+17, 1.313813777326696e+17, 1.313813777418883e+17, 1.31381377746732e+17, 1.31381377749857e+17, 1.313813777612632e+17, 1.31381377769232e+17, 1.313813777762632e+17, 1.313813777834508e+17, 1.313813777915758e+17, 1.313813777993883e+17, 1.313813778050132e+17, 1.313813778122008e+17, 1.313813778222007e+17, 1.313813778247008e+17, 1.313813778270445e+17, 1.31381377839232e+17, 1.313813778425133e+17, 1.313813778481382e+17, 1.313813778534508e+17, 1.313813778607945e+17, 1.313813778678257e+17, 1.313813778703258e+17, 1.313813778822008e+17, 1.313813778847008e+17, 1.313813778934508e+17, 1.313813779025133e+17, 1.313813779059508e+17, 1.313813779122007e+17, 1.313813779193883e+17, 1.31381377926107e+17, 1.313813779331383e+17, 1.313813779395444e+17, 1.313813779478258e+17, 1.313813779518883e+17, 1.313813779590757e+17, 1.31381377966107e+17, 1.313813779732945e+17, 1.313813779803258e+17, 1.31381377987982e+17, 1.31381377997982e+17, 1.31381378003607e+17, 1.313813780107945e+17, 1.313813780178257e+17, 1.313813780256383e+17, 1.313813780303258e+17, 1.313813780326694e+17, 1.313813780384508e+17, 1.31381378049232e+17, 1.313813780572008e+17, 1.313813780643884e+17, 1.313813780715758e+17, 1.313813780739195e+17, 1.313813780859507e+17, 1.31381378090482e+17, 1.31381378097982e+17, 1.313813781062633e+17, 1.313813781109507e+17, 1.31381378119232e+17, 1.313813781240758e+17, 1.313813781309508e+17, 1.313813781373571e+17, 1.313813781456383e+17, 1.313813781526694e+17, 1.31381378161732e+17, 1.313813781656381e+17, 1.313813781728257e+17, 1.313813781789196e+17, 1.31381378186107e+17, 1.313813781932945e+17, 1.313813782028257e+17, 1.313813782056383e+17, 1.313813782126696e+17, 1.313813782156383e+17, 1.31381378223607e+17, 1.31381378228607e+17, 1.313813782368883e+17, 1.313813782440758e+17, 1.313813782509508e+17, 1.313813782570445e+17, 1.313813782648571e+17, 1.313813782709508e+17, 1.313813782782945e+17, 1.313813782854821e+17, 1.31381378292357e+17, 1.313813783053257e+17, 1.313813783078257e+17, 1.313813783150132e+17, 1.313813783229819e+17, 1.31381378326732e+17, 1.313813783339195e+17, 1.313813783420445e+17, 1.313813783473569e+17, 1.313813783553258e+17, 1.313813783634508e+17, 1.313813783706383e+17, 1.313813783778258e+17, 1.313813783839195e+17, 1.313813783911069e+17, 1.313813783976695e+17, 1.313813784047008e+17, 1.313813784070445e+17, 1.313813784142321e+17, 1.313813784215758e+17, 1.313813784306383e+17, 1.313813784368883e+17, 1.313813784431382e+17, 1.313813784501696e+17, 1.313813784572008e+17, 1.313813784647008e+17, 1.313813784718883e+17, 1.313813784797007e+17, 1.313813784890758e+17, 1.31381378492357e+17, 1.313813784981384e+17, 1.31381378502357e+17, 1.313813785047007e+17, 1.31381378516732e+17, 1.313813785190757e+17, 1.313813785295444e+17, 1.313813785350132e+17, 1.313813785426696e+17, 1.313813785497007e+17, 1.313813785572008e+17, 1.313813785640758e+17, 1.313813785664195e+17, 1.313813785775132e+17, 1.313813785840756e+17, 1.313813785887633e+17, 1.313813785959508e+17, 1.31381378602982e+17, 1.313813786093883e+17, 1.313813786168882e+17, 1.31381378621732e+17, 1.313813786290757e+17, 1.313813786364195e+17, 1.31381378643607e+17, 1.313813786518883e+17, 1.313813786590757e+17, 1.313813786618883e+17, 1.313813786742321e+17, 1.313813786806382e+17, 1.313813786878258e+17, 1.313813786951695e+17, 1.313813787020444e+17, 1.31381378708607e+17, 1.313813787168883e+17, 1.313813787250132e+17, 1.31381378732357e+17, 1.313813787395444e+17, 1.313813787468883e+17, 1.313813787542319e+17, 1.31381378762357e+17, 1.313813787697007e+17, 1.31381378777982e+17, 1.31381378786107e+17, 1.313813787942321e+17, 1.31381378799857e+17, 1.313813788059507e+17, 1.313813788131382e+17, 1.313813788200132e+17, 1.313813788265757e+17, 1.313813788339195e+17, 1.313813788411069e+17, 1.313813788481382e+17, 1.31381378854857e+17, 1.313813788572008e+17, 1.31381378869857e+17, 1.313813788722007e+17, 1.313813788801695e+17, 1.313813788856383e+17, 1.313813788928257e+17, 1.313813789000132e+17, 1.313813789072008e+17, 1.313813789143884e+17, 1.313813789217321e+17, 1.31381378932982e+17, 1.31381378935482e+17, 1.313813789434508e+17, 1.313813789487633e+17, 1.31381378956732e+17, 1.313813789640758e+17, 1.313813789722007e+17, 1.31381378978607e+17, 1.313813789857944e+17, 1.313813789940758e+17, 1.313813790025133e+17, 1.31381379008607e+17, 1.313813790159507e+17, 1.31381379022982e+17, 1.313813790293883e+17, 1.313813790365757e+17, 1.313813790465757e+17, 1.313813790503258e+17, 1.31381379059857e+17, 1.313813790631383e+17, 1.313813790709508e+17, 1.313813790784508e+17, 1.313813790857946e+17, 1.313813790918883e+17, 1.313813790942321e+17, 1.313813791073569e+17, 1.313813791145445e+17, 1.313813791226696e+17, 1.313813791326696e+17, 1.313813791381382e+17, 1.313813791468883e+17, 1.313813791514195e+17, 1.31381379159857e+17, 1.313813791672008e+17, 1.313813791743884e+17, 1.313813791820444e+17, 1.313813791882945e+17, 1.313813791982944e+17, 1.31381379203607e+17, 1.313813792107945e+17, 1.313813792178257e+17, 1.313813792243882e+17, 1.313813792307945e+17, 1.313813792411071e+17, 1.313813792453258e+17, 1.313813792514195e+17, 1.313813792537632e+17, 1.313813792647008e+17, 1.31381379276107e+17, 1.313813792784507e+17, 1.31381379286732e+17, 1.31381379291732e+17, 1.313813793022007e+17, 1.313813793075132e+17, 1.31381379309857e+17, 1.313813793220445e+17, 1.313813793243884e+17, 1.313813793342321e+17, 1.313813793365757e+17, 1.313813793489194e+17, 1.313813793528257e+17, 1.313813793562632e+17, 1.313813793670445e+17, 1.313813793745445e+17, 1.313813793809508e+17, 1.31381379387982e+17, 1.313813793953257e+17, 1.313813794039196e+17, 1.313813794109507e+17, 1.313813794181382e+17, 1.313813794251695e+17, 1.313813794312632e+17, 1.313813794384507e+17, 1.313813794457946e+17, 1.313813794528257e+17, 1.31381379460482e+17, 1.313813794665757e+17, 1.31381379478607e+17, 1.313813794817321e+17, 1.313813794887633e+17, 1.313813794976695e+17, 1.31381379502982e+17, 1.313813795114195e+17, 1.313813795187633e+17, 1.313813795256383e+17, 1.31381379532357e+17, 1.313813795407945e+17, 1.313813795478258e+17, 1.31381379556107e+17, 1.313813795609508e+17, 1.313813795665757e+17, 1.313813795739195e+17, 1.313813795768882e+17, 1.313813795818883e+17, 1.313813795934508e+17, 1.313813796004819e+17, 1.313813796079821e+17, 1.31381379616107e+17, 1.313813796259507e+17, 1.313813796284507e+17, 1.313813796307945e+17, 1.313813796412632e+17, 1.313813796453257e+17, 1.31381379652982e+17, 1.313813796603258e+17, 1.313813796672008e+17, 1.313813796753257e+17, 1.313813796825133e+17, 1.31381379689857e+17, 1.313813796982945e+17, 1.313813797045445e+17, 1.313813797128257e+17, 1.313813797248571e+17, 1.313813797281382e+17, 1.313813797343884e+17, 1.313813797389196e+17, 1.313813797473571e+17, 1.313813797526696e+17, 1.313813797617321e+17, 1.313813797645444e+17, 1.313813797739196e+17, 1.31381379776732e+17, 1.313813797828257e+17, 1.313813797875132e+17, 1.313813797943882e+17, 1.313813798014195e+17, 1.313813798039195e+17, 1.313813798151695e+17, 1.31381379817982e+17, 1.31381379826107e+17, 1.313813798342321e+17, 1.31381379841732e+17, 1.313813798490757e+17, 1.313813798553257e+17, 1.313813798626696e+17, 1.313813798687633e+17, 1.313813798756383e+17, 1.313813798834508e+17, 1.313813798903256e+17, 1.313813798981382e+17, 1.31381379905482e+17, 1.313813799120445e+17, 1.313813799228257e+17, 1.31381379926107e+17, 1.313813799345445e+17, 1.313813799425133e+17, 1.313813799472008e+17, 1.313813799543884e+17, 1.313813799626694e+17, 1.313813799700132e+17, 1.313813799772006e+17, 1.313813799853258e+17, 1.31381379991732e+17, 1.313813799989196e+17, 1.313813800059508e+17, 1.31381380012982e+17, 1.31381380022357e+17, 1.313813800273571e+17, 1.313813800378258e+17, 1.31381380042982e+17, 1.313813800503258e+17, 1.313813800573569e+17, 1.313813800604819e+17, 1.313813800728257e+17, 1.313813800793883e+17, 1.313813800865756e+17, 1.31381380093607e+17, 1.313813800965757e+17, 1.313813801089196e+17, 1.313813801147008e+17, 1.313813801222007e+17, 1.313813801245445e+17, 1.313813801365757e+17, 1.313813801442319e+17, 1.313813801497007e+17, 1.313813801565757e+17, 1.313813801647008e+17, 1.313813801704819e+17, 1.313813801814195e+17, 1.313813801839195e+17, 1.313813801920444e+17, 1.313813801956383e+17, 1.313813802028257e+17, 1.313813802093883e+17, 1.313813802151695e+17, 1.31381380222357e+17, 1.313813802297007e+17, 1.313813802406382e+17, 1.313813802448571e+17, 1.313813802522008e+17, 1.313813802550132e+17, 1.313813802673571e+17, 1.313813802720445e+17, 1.313813802828257e+17, 1.313813802851694e+17, 1.313813802875132e+17, 1.313813802976695e+17, 1.31381380302982e+17, 1.313813803095444e+17, 1.313813803176695e+17, 1.313813803201695e+17, 1.313813803320444e+17, 1.313813803343882e+17, 1.313813803440758e+17, 1.313813803464195e+17, 1.313813803557946e+17, 1.313813803600132e+17, 1.313813803668883e+17, 1.313813803732945e+17, 1.313813803814195e+17, 1.313813803887633e+17, 1.313813803912632e+17, 1.313813804032946e+17, 1.31381380409857e+17, 1.313813804182944e+17, 1.313813804245445e+17, 1.313813804315757e+17, 1.313813804339195e+17, 1.313813804462632e+17, 1.313813804547007e+17, 1.313813804586071e+17, 1.313813804665757e+17, 1.313813804747007e+17, 1.313813804817321e+17, 1.313813804889196e+17, 1.313813804970445e+17, 1.313813805045444e+17, 1.313813805093883e+17, 1.313813805164195e+17, 1.313813805234508e+17, 1.313813805306382e+17, 1.31381380537982e+17, 1.313813805437633e+17, 1.313813805515758e+17, 1.31381380558607e+17, 1.313813805611069e+17, 1.31381380572982e+17, 1.313813805753258e+17, 1.313813805851695e+17, 1.31381380589232e+17, 1.313813805917321e+17, 1.313813806039195e+17, 1.313813806120444e+17, 1.313813806175132e+17, 1.313813806240756e+17, 1.313813806314195e+17, 1.313813806389196e+17, 1.313813806465757e+17, 1.313813806537633e+17, 1.313813806611071e+17, 1.313813806672008e+17, 1.313813806745445e+17, 1.313813806818883e+17, 1.313813806842321e+17, 1.313813806964195e+17, 1.313813807026694e+17, 1.313813807109508e+17, 1.313813807182944e+17, 1.313813807251695e+17, 1.313813807315757e+17, 1.313813807387633e+17, 1.313813807487631e+17, 1.313813807539195e+17, 1.313813807614195e+17, 1.31381380768607e+17, 1.313813807782945e+17, 1.313813807853258e+17, 1.313813807909508e+17, 1.313813807982945e+17, 1.313813808070445e+17, 1.313813808118883e+17, 1.313813808218883e+17, 1.313813808272008e+17, 1.313813808343882e+17, 1.313813808437633e+17, 1.313813808484507e+17, 1.313813808553257e+17, 1.31381380862357e+17, 1.313813808707945e+17, 1.313813808742321e+17, 1.31381380882982e+17, 1.313813808868883e+17, 1.313813808942321e+17, 1.313813809011069e+17, 1.313813809082945e+17, 1.313813809106382e+17, 1.313813809225132e+17, 1.31381380924857e+17, 1.313813809337632e+17, 1.313813809401695e+17, 1.313813809482945e+17, 1.313813809531383e+17, 1.313813809603258e+17, 1.31381380969232e+17},
			             {1.31381364866107e+17, 1.313813648847008e+17},
			             {1.313813786878258e+17, 1.31381378708607e+17},
			             {1.31381380969232e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}}, {{}, {}}, {{}};
		}
	}
}
