netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 18;
			channels = 6;
			categories = 75;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0,  50.0,  15.0,  15.0,  15.0,  15.0,  15.0, 172.4, 181.1, 178.8, 186.6, 179.3, 130.3, 120.1, 112.4, 107.0, 102.6,  99.1;
			max_depth =  70.4, 173.3, 250.9, 185.1, 244.7, 223.7, 206.6, 197.8, 189.2, 185.6, 198.6, 185.7, 205.7, 152.7, 144.6, 166.3, 153.0, 146.4;
			start_time = 127767684100681984, 127767684100681984, 127767699080681984, 127767684410681984, 127767694480681984, 127767691460681984, 127767687110681984, 127767706080681984, 127767702330681984, 127767702600681984, 127767703200681984, 127767703100681984, 127767707040681984, 127767691700681984, 127767692400681984, 127767693370681984, 127767691610681984, 127767688240681984;
			end_time = 127767684410681984, 127767684410681984, 127767718339432064, 127767687110681984, 127767699080681984, 127767694480681984, 127767691460681984, 127767706210681984, 127767702430681984, 127767702640681984, 127767703240681984, 127767703160681984, 127767718339432064, 127767692170681984, 127767692610681984, 127767693630681984, 127767692370681984, 127767689900681984;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "6", "5014", "6", "6", "6", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "12", "12", "12", "12", "12", "12", "12", "12", "12", "12", "12", "12";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 0.4, 0.6, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 74, 75;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "364";
			region_channels = 63, 63, 63, 63, 63, 63, 63,  0, 16, 16, 16, 16, 16, 63, 63, 63, 63, 63;
			mask_times = {1.27767684100682e+17, 1.27767684110682e+17, 1.27767684120682e+17, 1.27767684130682e+17, 1.27767684140682e+17, 1.27767684150682e+17, 1.27767684160682e+17, 1.27767684170682e+17, 1.27767684180682e+17, 1.27767684190682e+17, 1.27767684200682e+17, 1.27767684210682e+17, 1.27767684220682e+17, 1.27767684230682e+17, 1.27767684240682e+17, 1.27767684250682e+17, 1.27767684260682e+17, 1.27767684270682e+17, 1.27767684280682e+17, 1.27767684290682e+17, 1.27767684300682e+17, 1.27767684310682e+17, 1.27767684320682e+17, 1.27767684330682e+17, 1.27767684340682e+17, 1.27767684350682e+17, 1.27767684360682e+17, 1.27767684370682e+17, 1.27767684380682e+17, 1.27767684390682e+17, 1.27767684400682e+17, 1.27767684410682e+17},
			             {1.27767684100682e+17, 1.27767684110682e+17, 1.27767684120682e+17, 1.27767684130682e+17, 1.27767684140682e+17, 1.27767684150682e+17, 1.27767684160682e+17, 1.27767684170682e+17, 1.27767684180682e+17, 1.27767684190682e+17, 1.27767684200682e+17, 1.27767684210682e+17, 1.27767684220682e+17, 1.27767684230682e+17, 1.27767684240682e+17, 1.27767684250682e+17, 1.27767684260682e+17, 1.27767684270682e+17, 1.27767684280682e+17, 1.27767684290682e+17, 1.27767684300682e+17, 1.27767684310682e+17, 1.27767684320682e+17, 1.27767684330682e+17, 1.27767684340682e+17, 1.27767684350682e+17, 1.27767684360682e+17, 1.27767684370682e+17, 1.27767684380682e+17, 1.27767684390682e+17, 1.27767684400682e+17, 1.27767684410682e+17},
			             {1.27767699080682e+17, 1.27767699090682e+17, 1.27767699100682e+17, 1.27767699110682e+17, 1.27767699120682e+17, 1.277676991306821e+17, 1.27767699140682e+17, 1.27767699150682e+17, 1.27767699160682e+17, 1.27767699170682e+17, 1.27767699180682e+17, 1.27767699190682e+17, 1.27767699200682e+17, 1.27767699210682e+17, 1.27767699220682e+17, 1.27767699230682e+17, 1.27767699240682e+17, 1.27767699250682e+17, 1.27767699260682e+17, 1.27767699270682e+17, 1.27767699280682e+17, 1.27767699290682e+17, 1.27767699300682e+17, 1.27767699310682e+17, 1.27767699320682e+17, 1.27767699330682e+17, 1.27767699340682e+17, 1.27767699350682e+17, 1.27767699360682e+17, 1.27767699370682e+17, 1.27767699380682e+17, 1.277676993906821e+17, 1.27767699400682e+17, 1.27767699410682e+17, 1.27767699420682e+17, 1.27767699430682e+17, 1.27767699440682e+17, 1.27767699450682e+17, 1.27767699460682e+17, 1.27767699470682e+17, 1.27767699480682e+17, 1.27767699490682e+17, 1.27767699500682e+17, 1.27767699510682e+17, 1.27767699520682e+17, 1.27767699530682e+17, 1.27767699540682e+17, 1.27767699550682e+17, 1.27767699560682e+17, 1.27767699570682e+17, 1.27767699580682e+17, 1.27767699590682e+17, 1.27767699600682e+17, 1.27767699610682e+17, 1.27767699620682e+17, 1.27767699630682e+17, 1.27767699640682e+17, 1.27767699650682e+17, 1.27767699660682e+17, 1.27767699670682e+17, 1.27767699680682e+17, 1.27767699690682e+17, 1.27767699700682e+17, 1.27767699710682e+17, 1.27767699720682e+17, 1.27767699730682e+17, 1.27767699740682e+17, 1.27767699750682e+17, 1.277676997606821e+17, 1.27767699770682e+17, 1.27767699780682e+17, 1.27767699790682e+17, 1.27767699800682e+17, 1.27767699810682e+17, 1.27767699820682e+17, 1.27767699830682e+17, 1.27767699840682e+17, 1.27767699850682e+17, 1.27767699860682e+17, 1.27767699870682e+17, 1.27767699880682e+17, 1.27767699890682e+17, 1.27767699900682e+17, 1.27767699910682e+17, 1.27767699920682e+17, 1.27767699930682e+17, 1.27767699940682e+17, 1.27767699950682e+17, 1.27767699960682e+17, 1.27767699970682e+17, 1.27767699980682e+17, 1.27767699990682e+17, 1.27767700000682e+17, 1.27767700010682e+17, 1.277677000206821e+17, 1.27767700030682e+17, 1.27767700040682e+17, 1.27767700050682e+17, 1.27767700060682e+17, 1.27767700070682e+17, 1.27767700080682e+17, 1.27767700090682e+17, 1.27767700100682e+17, 1.27767700110682e+17, 1.27767700120682e+17, 1.27767700130682e+17, 1.27767700140682e+17, 1.27767700150682e+17, 1.27767700160682e+17, 1.27767700170682e+17, 1.27767700180682e+17, 1.27767700190682e+17, 1.27767700200682e+17, 1.27767700210682e+17, 1.27767700220682e+17, 1.27767700230682e+17, 1.27767700240682e+17, 1.27767700250682e+17, 1.27767700260682e+17, 1.27767700270682e+17, 1.277677002806821e+17, 1.27767700290682e+17, 1.27767700300682e+17, 1.27767700310682e+17, 1.27767700320682e+17, 1.27767700330682e+17, 1.27767700340682e+17, 1.27767700350682e+17, 1.27767700360682e+17, 1.27767700370682e+17, 1.27767700380682e+17, 1.27767700390682e+17, 1.27767700400682e+17, 1.27767700410682e+17, 1.27767700420682e+17, 1.27767700430682e+17, 1.27767700440682e+17, 1.27767700450682e+17, 1.277677004608383e+17, 1.27767700470682e+17, 1.27767700480682e+17, 1.27767700490682e+17, 1.27767700500682e+17, 1.27767700510682e+17, 1.27767700520682e+17, 1.27767700530682e+17, 1.27767700540682e+17, 1.27767700550682e+17, 1.27767700560682e+17, 1.27767700570682e+17, 1.27767700580682e+17, 1.27767700590682e+17, 1.27767700600682e+17, 1.27767700610682e+17, 1.27767700620682e+17, 1.27767700630682e+17, 1.27767700640682e+17, 1.27767700650682e+17, 1.27767700660682e+17, 1.27767700670682e+17, 1.27767700680682e+17, 1.27767700690682e+17, 1.27767700700682e+17, 1.27767700710682e+17, 1.27767700720682e+17, 1.27767700730682e+17, 1.27767700740682e+17, 1.27767700750682e+17, 1.27767700760682e+17, 1.27767700770682e+17, 1.27767700780682e+17, 1.27767700790682e+17, 1.27767700800682e+17, 1.27767700810682e+17, 1.27767700820682e+17, 1.27767700830682e+17, 1.27767700840682e+17, 1.27767700850682e+17, 1.27767700860682e+17, 1.27767700870682e+17, 1.27767700880682e+17, 1.27767700890682e+17, 1.27767700900682e+17, 1.277677009106821e+17, 1.27767700920682e+17, 1.27767700930682e+17, 1.27767700940682e+17, 1.27767700950682e+17, 1.27767700960682e+17, 1.27767700970682e+17, 1.27767700980682e+17, 1.27767700990682e+17, 1.27767701000682e+17, 1.27767701010682e+17, 1.27767701020682e+17, 1.27767701030682e+17, 1.27767701040682e+17, 1.27767701050682e+17, 1.27767701060682e+17, 1.27767701070682e+17, 1.27767701080682e+17, 1.27767701090682e+17, 1.27767701100682e+17, 1.27767701110682e+17, 1.27767701120682e+17, 1.27767701130682e+17, 1.27767701140682e+17, 1.27767701150682e+17, 1.27767701160682e+17, 1.277677011706821e+17, 1.27767701180682e+17, 1.27767701190682e+17, 1.27767701200682e+17, 1.27767701210682e+17, 1.27767701220682e+17, 1.27767701230682e+17, 1.27767701240682e+17, 1.27767701250682e+17, 1.27767701260682e+17, 1.27767701270682e+17, 1.27767701280682e+17, 1.27767701290682e+17, 1.27767701300682e+17, 1.27767701310682e+17, 1.27767701320682e+17, 1.27767701330682e+17, 1.27767701340682e+17, 1.27767701350682e+17, 1.27767701360682e+17, 1.27767701370682e+17, 1.27767701380682e+17, 1.27767701390682e+17, 1.27767701400682e+17, 1.27767701410682e+17, 1.27767701420682e+17, 1.277677014306821e+17, 1.27767701440682e+17, 1.27767701450682e+17, 1.27767701460682e+17, 1.27767701470682e+17, 1.27767701480682e+17, 1.27767701490682e+17, 1.27767701500682e+17, 1.27767701510682e+17, 1.27767701520682e+17, 1.27767701530682e+17, 1.27767701540682e+17, 1.27767701550682e+17, 1.27767701560682e+17, 1.27767701570682e+17, 1.27767701580682e+17, 1.27767701590682e+17, 1.27767701600682e+17, 1.27767701610682e+17, 1.27767701620682e+17, 1.27767701630682e+17, 1.27767701640682e+17, 1.27767701650682e+17, 1.27767701660682e+17, 1.27767701670682e+17, 1.27767701680682e+17, 1.27767701690682e+17, 1.27767701700682e+17, 1.27767701710682e+17, 1.27767701720682e+17, 1.27767701730682e+17, 1.27767701740682e+17, 1.27767701750682e+17, 1.27767701760682e+17, 1.27767701770682e+17, 1.27767701780682e+17, 1.27767701790682e+17, 1.277677018006821e+17, 1.27767701810682e+17, 1.27767701820682e+17, 1.27767701830682e+17, 1.27767701840682e+17, 1.27767701850682e+17, 1.27767701860682e+17, 1.27767701870682e+17, 1.27767701880682e+17, 1.27767701890682e+17, 1.27767701900682e+17, 1.27767701910682e+17, 1.27767701920682e+17, 1.27767701930682e+17, 1.27767701940682e+17, 1.27767701950682e+17, 1.27767701960682e+17, 1.27767701970682e+17, 1.27767701980682e+17, 1.27767701990682e+17, 1.27767702000682e+17, 1.27767702010682e+17, 1.27767702020682e+17, 1.27767702030682e+17, 1.27767702040682e+17, 1.27767702050682e+17, 1.277677020606821e+17, 1.27767702070682e+17, 1.27767702080682e+17, 1.27767702090682e+17, 1.27767702100682e+17, 1.27767702110682e+17, 1.27767702120682e+17, 1.27767702130682e+17, 1.27767702140682e+17, 1.27767702150682e+17, 1.27767702160682e+17, 1.27767702170682e+17, 1.27767702180682e+17, 1.27767702190682e+17, 1.27767702200682e+17, 1.27767702210682e+17, 1.27767702220682e+17, 1.27767702230682e+17, 1.27767702240682e+17, 1.27767702250682e+17, 1.27767702260682e+17, 1.27767702270682e+17, 1.27767702280682e+17, 1.27767702290682e+17, 1.27767702300682e+17, 1.27767702310682e+17, 1.277677023206821e+17, 1.27767702330682e+17, 1.27767702340682e+17, 1.27767702350682e+17, 1.27767702360682e+17, 1.27767702370682e+17, 1.27767702380682e+17, 1.27767702390682e+17, 1.27767702400682e+17, 1.27767702410682e+17, 1.27767702420682e+17, 1.27767702430682e+17, 1.27767702440682e+17, 1.27767702450682e+17, 1.27767702460682e+17, 1.27767702470682e+17, 1.27767702480682e+17, 1.27767702490682e+17, 1.27767702500682e+17, 1.27767702510682e+17, 1.27767702520682e+17, 1.27767702530682e+17, 1.27767702540682e+17, 1.27767702550682e+17, 1.27767702560682e+17, 1.27767702570682e+17, 1.27767702580682e+17, 1.27767702590682e+17, 1.27767702600682e+17, 1.27767702610682e+17, 1.27767702620682e+17, 1.27767702630682e+17, 1.27767702640682e+17, 1.27767702650682e+17, 1.27767702660682e+17, 1.27767702670682e+17, 1.27767702680682e+17, 1.277677026906821e+17, 1.27767702700682e+17, 1.27767702710682e+17, 1.27767702720682e+17, 1.27767702730682e+17, 1.27767702740682e+17, 1.27767702750682e+17, 1.27767702760682e+17, 1.27767702770682e+17, 1.27767702780682e+17, 1.27767702790682e+17, 1.27767702800682e+17, 1.27767702810682e+17, 1.27767702820682e+17, 1.27767702830682e+17, 1.27767702840682e+17, 1.27767702850682e+17, 1.27767702860682e+17, 1.27767702870682e+17, 1.27767702880682e+17, 1.27767702890682e+17, 1.27767702900682e+17, 1.27767702910682e+17, 1.27767702920682e+17, 1.27767702930682e+17, 1.27767702940682e+17, 1.277677029506821e+17, 1.27767702960682e+17, 1.27767702970682e+17, 1.27767702980682e+17, 1.27767702990682e+17, 1.27767703000682e+17, 1.27767703010682e+17, 1.27767703020682e+17, 1.27767703030682e+17, 1.27767703040682e+17, 1.27767703050682e+17, 1.27767703060682e+17, 1.27767703070682e+17, 1.27767703080682e+17, 1.27767703090682e+17, 1.27767703100682e+17, 1.27767703110682e+17, 1.27767703120682e+17, 1.27767703130682e+17, 1.27767703140682e+17, 1.27767703150682e+17, 1.27767703160682e+17, 1.27767703170682e+17, 1.27767703180682e+17, 1.27767703190682e+17, 1.27767703200682e+17, 1.277677032106821e+17, 1.27767703220682e+17, 1.27767703230682e+17, 1.27767703240682e+17, 1.27767703250682e+17, 1.27767703260682e+17, 1.27767703270682e+17, 1.27767703280682e+17, 1.27767703290682e+17, 1.27767703300682e+17, 1.27767703310682e+17, 1.27767703320682e+17, 1.27767703330682e+17, 1.27767703340682e+17, 1.27767703350682e+17, 1.27767703360682e+17, 1.27767703370682e+17, 1.27767703380682e+17, 1.27767703390682e+17, 1.27767703400682e+17, 1.27767703410682e+17, 1.27767703420682e+17, 1.27767703430682e+17, 1.27767703440682e+17, 1.27767703450682e+17, 1.27767703460682e+17, 1.27767703470682e+17, 1.27767703480682e+17, 1.27767703490682e+17, 1.27767703500682e+17, 1.27767703510682e+17, 1.27767703520682e+17, 1.27767703530682e+17, 1.27767703540682e+17, 1.27767703550682e+17, 1.27767703560682e+17, 1.27767703570682e+17, 1.277677035806821e+17, 1.27767703590682e+17, 1.27767703600682e+17, 1.27767703610682e+17, 1.27767703620682e+17, 1.27767703630682e+17, 1.27767703640682e+17, 1.27767703650682e+17, 1.27767703660682e+17, 1.27767703670682e+17, 1.27767703680682e+17, 1.27767703690682e+17, 1.27767703700682e+17, 1.27767703710682e+17, 1.27767703720682e+17, 1.27767703730682e+17, 1.27767703740682e+17, 1.27767703750682e+17, 1.27767703760682e+17, 1.27767703770682e+17, 1.27767703780682e+17, 1.27767703790682e+17, 1.27767703800682e+17, 1.27767703810682e+17, 1.27767703820682e+17, 1.27767703830682e+17, 1.277677038406821e+17, 1.27767703850682e+17, 1.27767703860682e+17, 1.27767703870682e+17, 1.27767703880682e+17, 1.27767703890682e+17, 1.27767703900682e+17, 1.27767703910682e+17, 1.27767703920682e+17, 1.27767703930682e+17, 1.27767703940682e+17, 1.27767703950682e+17, 1.27767703960682e+17, 1.27767703970682e+17, 1.27767703980682e+17, 1.27767703990682e+17, 1.27767704000682e+17, 1.27767704010682e+17, 1.27767704020682e+17, 1.27767704030682e+17, 1.27767704040682e+17, 1.27767704050682e+17, 1.27767704060682e+17, 1.27767704070682e+17, 1.27767704080682e+17, 1.27767704090682e+17, 1.277677041006821e+17, 1.27767704110682e+17, 1.27767704120682e+17, 1.27767704130682e+17, 1.27767704140682e+17, 1.27767704150682e+17, 1.27767704160682e+17, 1.27767704170682e+17, 1.27767704180682e+17, 1.27767704190682e+17, 1.27767704200682e+17, 1.27767704210682e+17, 1.27767704220682e+17, 1.27767704230682e+17, 1.27767704240682e+17, 1.27767704250682e+17, 1.27767704260682e+17, 1.27767704270682e+17, 1.27767704280682e+17, 1.27767704290682e+17, 1.27767704300682e+17, 1.27767704310682e+17, 1.27767704320682e+17, 1.27767704330682e+17, 1.27767704340682e+17, 1.27767704350682e+17, 1.27767704360682e+17, 1.27767704370682e+17, 1.27767704380682e+17, 1.27767704390682e+17, 1.27767704400682e+17, 1.27767704410682e+17, 1.27767704420682e+17, 1.27767704430682e+17, 1.27767704440682e+17, 1.27767704450682e+17, 1.27767704460682e+17, 1.27767704470682e+17, 1.27767704480682e+17, 1.27767704490682e+17, 1.27767704500682e+17, 1.27767704510682e+17, 1.27767704520682e+17, 1.27767704530682e+17, 1.27767704540682e+17, 1.27767704550682e+17, 1.27767704560682e+17, 1.27767704570682e+17, 1.27767704580682e+17, 1.27767704590682e+17, 1.27767704600682e+17, 1.27767704610682e+17, 1.27767704620682e+17, 1.27767704630682e+17, 1.27767704640682e+17, 1.27767704650682e+17, 1.27767704660682e+17, 1.27767704670682e+17, 1.27767704680682e+17, 1.27767704690682e+17, 1.27767704700682e+17, 1.27767704710682e+17, 1.27767704720682e+17, 1.277677047306821e+17, 1.27767704740682e+17, 1.27767704750682e+17, 1.27767704760682e+17, 1.27767704770682e+17, 1.27767704780682e+17, 1.27767704790682e+17, 1.27767704800682e+17, 1.27767704810682e+17, 1.27767704820682e+17, 1.27767704830682e+17, 1.27767704840682e+17, 1.27767704850682e+17, 1.27767704860682e+17, 1.27767704870682e+17, 1.27767704880682e+17, 1.27767704890682e+17, 1.27767704900682e+17, 1.27767704910682e+17, 1.27767704920682e+17, 1.27767704930682e+17, 1.27767704940682e+17, 1.27767704950682e+17, 1.27767704960682e+17, 1.27767704970682e+17, 1.27767704980682e+17, 1.277677049906821e+17, 1.27767705000682e+17, 1.27767705010682e+17, 1.27767705020682e+17, 1.27767705030682e+17, 1.27767705040682e+17, 1.27767705050682e+17, 1.27767705060682e+17, 1.27767705070682e+17, 1.27767705080682e+17, 1.27767705090682e+17, 1.27767705100682e+17, 1.27767705110682e+17, 1.27767705120682e+17, 1.27767705130682e+17, 1.27767705140682e+17, 1.27767705150682e+17, 1.27767705160682e+17, 1.27767705170682e+17, 1.27767705180682e+17, 1.27767705190682e+17, 1.27767705200682e+17, 1.27767705210682e+17, 1.27767705220682e+17, 1.27767705230682e+17, 1.27767705240682e+17, 1.277677052506821e+17, 1.27767705260682e+17, 1.27767705270682e+17, 1.27767705280682e+17, 1.27767705290682e+17, 1.27767705300682e+17, 1.27767705310682e+17, 1.27767705320682e+17, 1.27767705330682e+17, 1.27767705340682e+17, 1.27767705350682e+17, 1.27767705360682e+17, 1.27767705370682e+17, 1.27767705380682e+17, 1.27767705390682e+17, 1.27767705400682e+17, 1.27767705410682e+17, 1.27767705420682e+17, 1.27767705430682e+17, 1.27767705440682e+17, 1.27767705450682e+17, 1.27767705460682e+17, 1.27767705470682e+17, 1.27767705480682e+17, 1.27767705490682e+17, 1.27767705500682e+17, 1.27767705510682e+17, 1.27767705520682e+17, 1.27767705530682e+17, 1.27767705540682e+17, 1.27767705550682e+17, 1.27767705560682e+17, 1.27767705570682e+17, 1.27767705580682e+17, 1.27767705590682e+17, 1.27767705600682e+17, 1.27767705610682e+17, 1.277677056206821e+17, 1.27767705630682e+17, 1.27767705640682e+17, 1.27767705650682e+17, 1.27767705660682e+17, 1.27767705670682e+17, 1.27767705680682e+17, 1.27767705690682e+17, 1.27767705700682e+17, 1.27767705710682e+17, 1.27767705720682e+17, 1.27767705730682e+17, 1.27767705740682e+17, 1.27767705750682e+17, 1.27767705760682e+17, 1.27767705770682e+17, 1.27767705780682e+17, 1.27767705790682e+17, 1.27767705800682e+17, 1.27767705810682e+17, 1.27767705820682e+17, 1.27767705830682e+17, 1.27767705840682e+17, 1.27767705850682e+17, 1.27767705860682e+17, 1.27767705870682e+17, 1.277677058806821e+17, 1.27767705890682e+17, 1.27767705900682e+17, 1.27767705910682e+17, 1.27767705920682e+17, 1.27767705930682e+17, 1.27767705940682e+17, 1.27767705950682e+17, 1.27767705960682e+17, 1.27767705970682e+17, 1.27767705980682e+17, 1.27767705990682e+17, 1.27767706000682e+17, 1.27767706010682e+17, 1.27767706020682e+17, 1.27767706030682e+17, 1.27767706040682e+17, 1.27767706050682e+17, 1.27767706060682e+17, 1.27767706070682e+17, 1.27767706080682e+17, 1.27767706090682e+17, 1.27767706100682e+17, 1.27767706110682e+17, 1.27767706120682e+17, 1.27767706130682e+17, 1.277677061406821e+17, 1.27767706150682e+17, 1.27767706160682e+17, 1.27767706170682e+17, 1.27767706180682e+17, 1.27767706190682e+17, 1.27767706200682e+17, 1.27767706210682e+17, 1.27767706220682e+17, 1.27767706230682e+17, 1.27767706240682e+17, 1.27767706250682e+17, 1.27767706260682e+17, 1.27767706270682e+17, 1.27767706280682e+17, 1.27767706290682e+17, 1.27767706300682e+17, 1.27767706310682e+17, 1.27767706320682e+17, 1.27767706330682e+17, 1.27767706340682e+17, 1.27767706350682e+17, 1.27767706360682e+17, 1.27767706370682e+17, 1.27767706380682e+17, 1.27767706390682e+17, 1.27767706400682e+17, 1.27767706410682e+17, 1.27767706420682e+17, 1.27767706430682e+17, 1.27767706440682e+17, 1.27767706450682e+17, 1.27767706460682e+17, 1.27767706470682e+17, 1.27767706480682e+17, 1.27767706490682e+17, 1.27767706500682e+17, 1.277677065106821e+17, 1.27767706520682e+17, 1.27767706530682e+17, 1.27767706540682e+17, 1.27767706550682e+17, 1.27767706560682e+17, 1.27767706570682e+17, 1.27767706580682e+17, 1.27767706590682e+17, 1.27767706600682e+17, 1.27767706610682e+17, 1.27767706620682e+17, 1.27767706630682e+17, 1.27767706640682e+17, 1.27767706650682e+17, 1.27767706660682e+17, 1.27767706670682e+17, 1.27767706680682e+17, 1.27767706690682e+17, 1.27767706700682e+17, 1.27767706710682e+17, 1.27767706720682e+17, 1.27767706730682e+17, 1.27767706740682e+17, 1.27767706750682e+17, 1.27767706760682e+17, 1.277677067706821e+17, 1.27767706780682e+17, 1.27767706790682e+17, 1.27767706800682e+17, 1.27767706810682e+17, 1.27767706820682e+17, 1.27767706830682e+17, 1.27767706840682e+17, 1.27767706850682e+17, 1.27767706860682e+17, 1.27767706870682e+17, 1.27767706880682e+17, 1.27767706890682e+17, 1.27767706900682e+17, 1.27767706910682e+17, 1.27767706920682e+17, 1.27767706930682e+17, 1.27767706940682e+17, 1.27767706950682e+17, 1.27767706960682e+17, 1.27767706970682e+17, 1.27767706980682e+17, 1.27767706990682e+17, 1.27767707000682e+17, 1.27767707010682e+17, 1.27767707020682e+17, 1.277677070306821e+17, 1.27767707040682e+17, 1.27767707050682e+17, 1.27767707060682e+17, 1.27767707070682e+17, 1.27767707080682e+17, 1.27767707090682e+17, 1.27767707100682e+17, 1.27767707110682e+17, 1.27767707120682e+17, 1.27767707130682e+17, 1.27767707140682e+17, 1.27767707150682e+17, 1.27767707160682e+17, 1.27767707170682e+17, 1.27767707180682e+17, 1.27767707190682e+17, 1.27767707200682e+17, 1.27767707210682e+17, 1.27767707220682e+17, 1.27767707230682e+17, 1.27767707240682e+17, 1.27767707250682e+17, 1.27767707260682e+17, 1.27767707270682e+17, 1.27767707280682e+17, 1.27767707290682e+17, 1.27767707300682e+17, 1.27767707310682e+17, 1.27767707320682e+17, 1.27767707330682e+17, 1.27767707340682e+17, 1.27767707350682e+17, 1.27767707360682e+17, 1.27767707370682e+17, 1.27767707380682e+17, 1.27767707390682e+17, 1.27767707400682e+17, 1.27767707410682e+17, 1.27767707420682e+17, 1.27767707430682e+17, 1.27767707440682e+17, 1.27767707450682e+17, 1.27767707460682e+17, 1.27767707470682e+17, 1.27767707480682e+17, 1.27767707490682e+17, 1.27767707500682e+17, 1.27767707510682e+17, 1.27767707520682e+17, 1.27767707530682e+17, 1.27767707540682e+17, 1.27767707550682e+17, 1.27767707560682e+17, 1.27767707570682e+17, 1.27767707580682e+17, 1.27767707590682e+17, 1.27767707600682e+17, 1.27767707610682e+17, 1.27767707620682e+17, 1.27767707630682e+17, 1.27767707640682e+17, 1.27767707650682e+17, 1.277677076606821e+17, 1.27767707670682e+17, 1.27767707680682e+17, 1.27767707690682e+17, 1.27767707700682e+17, 1.27767707710682e+17, 1.27767707720682e+17, 1.27767707730682e+17, 1.27767707740682e+17, 1.27767707750682e+17, 1.27767707760682e+17, 1.27767707770682e+17, 1.27767707780682e+17, 1.27767707790682e+17, 1.27767707800682e+17, 1.27767707810682e+17, 1.27767707820682e+17, 1.27767707830682e+17, 1.27767707840682e+17, 1.27767707850682e+17, 1.27767707860682e+17, 1.27767707870682e+17, 1.27767707880682e+17, 1.27767707890682e+17, 1.27767707900682e+17, 1.27767707910682e+17, 1.277677079206821e+17, 1.27767707930682e+17, 1.27767707940682e+17, 1.27767707950682e+17, 1.27767707960682e+17, 1.27767707970682e+17, 1.27767707980682e+17, 1.27767707990682e+17, 1.27767708000682e+17, 1.27767708010682e+17, 1.27767708020682e+17, 1.27767708030682e+17, 1.27767708040682e+17, 1.27767708050682e+17, 1.27767708060682e+17, 1.27767708070682e+17, 1.27767708080682e+17, 1.27767708090682e+17, 1.27767708100682e+17, 1.27767708110682e+17, 1.27767708120682e+17, 1.27767708130682e+17, 1.27767708140682e+17, 1.27767708150682e+17, 1.27767708160682e+17, 1.27767708170682e+17, 1.277677081806821e+17, 1.27767708190682e+17, 1.27767708200682e+17, 1.27767708210682e+17, 1.27767708220682e+17, 1.27767708230682e+17, 1.27767708240682e+17, 1.27767708250682e+17, 1.27767708260682e+17, 1.27767708270682e+17, 1.27767708280682e+17, 1.27767708290682e+17, 1.27767708300682e+17, 1.27767708310682e+17, 1.27767708320682e+17, 1.27767708330682e+17, 1.27767708340682e+17, 1.27767708350682e+17, 1.27767708360682e+17, 1.27767708370682e+17, 1.27767708380682e+17, 1.27767708390682e+17, 1.27767708400682e+17, 1.27767708410682e+17, 1.27767708420682e+17, 1.27767708430682e+17, 1.27767708440682e+17, 1.27767708450682e+17, 1.27767708460682e+17, 1.27767708470682e+17, 1.27767708480682e+17, 1.27767708490682e+17, 1.27767708500682e+17, 1.27767708510682e+17, 1.27767708520682e+17, 1.27767708530682e+17, 1.27767708540682e+17, 1.277677085506821e+17, 1.27767708560682e+17, 1.27767708570682e+17, 1.27767708580682e+17, 1.27767708590682e+17, 1.27767708600682e+17, 1.27767708610682e+17, 1.27767708620682e+17, 1.27767708630682e+17, 1.27767708640682e+17, 1.27767708650682e+17, 1.27767708660682e+17, 1.27767708670682e+17, 1.27767708680682e+17, 1.27767708690682e+17, 1.27767708700682e+17, 1.27767708710682e+17, 1.27767708720682e+17, 1.27767708730682e+17, 1.27767708740682e+17, 1.27767708750682e+17, 1.27767708760682e+17, 1.27767708770682e+17, 1.27767708780682e+17, 1.27767708790682e+17, 1.27767708800682e+17, 1.277677088106821e+17, 1.27767708820682e+17, 1.27767708830682e+17, 1.27767708840682e+17, 1.27767708850682e+17, 1.27767708860682e+17, 1.27767708870682e+17, 1.27767708880682e+17, 1.27767708890682e+17, 1.27767708900682e+17, 1.27767708910682e+17, 1.27767708920682e+17, 1.27767708930682e+17, 1.27767708940682e+17, 1.27767708950682e+17, 1.27767708960682e+17, 1.27767708970682e+17, 1.27767708980682e+17, 1.27767708990682e+17, 1.27767709000682e+17, 1.27767709010682e+17, 1.27767709020682e+17, 1.27767709030682e+17, 1.27767709040682e+17, 1.27767709050682e+17, 1.27767709060682e+17, 1.277677090706821e+17, 1.27767709080682e+17, 1.27767709090682e+17, 1.27767709100682e+17, 1.27767709110682e+17, 1.27767709120682e+17, 1.27767709130682e+17, 1.27767709140682e+17, 1.27767709150682e+17, 1.27767709160682e+17, 1.27767709170682e+17, 1.27767709180682e+17, 1.27767709190682e+17, 1.27767709200682e+17, 1.27767709210682e+17, 1.27767709220682e+17, 1.27767709230682e+17, 1.27767709240682e+17, 1.27767709250682e+17, 1.27767709260682e+17, 1.27767709270682e+17, 1.27767709280682e+17, 1.27767709290682e+17, 1.27767709300682e+17, 1.27767709310682e+17, 1.27767709320682e+17, 1.27767709330682e+17, 1.27767709340682e+17, 1.27767709350682e+17, 1.27767709360682e+17, 1.27767709370682e+17, 1.27767709380682e+17, 1.27767709390682e+17, 1.27767709420682e+17, 1.27767709430682e+17, 1.277677094406821e+17, 1.27767709450682e+17, 1.27767709460682e+17, 1.27767709470682e+17, 1.27767709480682e+17, 1.27767709490682e+17, 1.27767709500682e+17, 1.27767709510682e+17, 1.27767709520682e+17, 1.27767709530682e+17, 1.27767709540682e+17, 1.27767709550682e+17, 1.27767709560682e+17, 1.27767709570682e+17, 1.27767709580682e+17, 1.27767709590682e+17, 1.27767709600682e+17, 1.27767709610682e+17, 1.27767709620682e+17, 1.27767709630682e+17, 1.27767709640682e+17, 1.27767709650682e+17, 1.27767709660682e+17, 1.27767709670682e+17, 1.27767709680682e+17, 1.27767709690682e+17, 1.277677097006821e+17, 1.27767709710682e+17, 1.27767709720682e+17, 1.27767709730682e+17, 1.27767709740682e+17, 1.27767709750682e+17, 1.27767709760682e+17, 1.27767709770682e+17, 1.27767709780682e+17, 1.27767709790682e+17, 1.27767709800682e+17, 1.27767709810682e+17, 1.27767709820682e+17, 1.27767709830682e+17, 1.27767709840682e+17, 1.27767709850682e+17, 1.27767709860682e+17, 1.27767709870682e+17, 1.27767709880682e+17, 1.27767709890682e+17, 1.27767709900682e+17, 1.27767709910682e+17, 1.27767709920682e+17, 1.27767709930682e+17, 1.27767709940682e+17, 1.27767709950682e+17, 1.277677099606821e+17, 1.27767709970682e+17, 1.27767709980682e+17, 1.27767709990682e+17, 1.27767710000682e+17, 1.27767710010682e+17, 1.27767710020682e+17, 1.27767710030682e+17, 1.27767710040682e+17, 1.27767710050682e+17, 1.27767710060682e+17, 1.27767710070682e+17, 1.27767710080682e+17, 1.27767710090682e+17, 1.27767710100682e+17, 1.27767710110682e+17, 1.27767710120682e+17, 1.27767710130682e+17, 1.27767710140682e+17, 1.27767710150682e+17, 1.27767710160682e+17, 1.27767710170682e+17, 1.27767710180682e+17, 1.27767710190682e+17, 1.27767710200682e+17, 1.27767710210682e+17, 1.27767710220682e+17, 1.27767710230682e+17, 1.27767710240682e+17, 1.27767710250682e+17, 1.27767710260682e+17, 1.27767710270682e+17, 1.27767710280682e+17, 1.27767710290682e+17, 1.27767710300682e+17, 1.27767710310682e+17, 1.27767710320682e+17, 1.277677103306821e+17, 1.27767710340682e+17, 1.27767710350682e+17, 1.27767710360682e+17, 1.27767710370682e+17, 1.27767710380682e+17, 1.27767710390682e+17, 1.27767710400682e+17, 1.27767710410682e+17, 1.27767710420682e+17, 1.27767710430682e+17, 1.27767710440682e+17, 1.27767710450682e+17, 1.27767710460682e+17, 1.27767710470682e+17, 1.27767710480682e+17, 1.27767710490682e+17, 1.27767710500682e+17, 1.27767710510682e+17, 1.27767710520682e+17, 1.27767710530682e+17, 1.27767710540682e+17, 1.27767710550682e+17, 1.27767710560682e+17, 1.27767710570682e+17, 1.27767710580682e+17, 1.277677105906821e+17, 1.27767710600682e+17, 1.27767710610682e+17, 1.27767710620682e+17, 1.27767710630682e+17, 1.27767710640682e+17, 1.27767710650682e+17, 1.27767710660682e+17, 1.27767710670682e+17, 1.27767710680682e+17, 1.27767710690682e+17, 1.27767710700682e+17, 1.27767710710682e+17, 1.27767710720682e+17, 1.27767710730682e+17, 1.27767710740682e+17, 1.27767710750682e+17, 1.27767710760682e+17, 1.27767710770682e+17, 1.27767710780682e+17, 1.27767710790682e+17, 1.27767710800682e+17, 1.27767710810682e+17, 1.27767710820682e+17, 1.27767710830682e+17, 1.27767710840682e+17, 1.277677108506821e+17, 1.27767710860682e+17, 1.277677108678696e+17, 1.27767710880682e+17, 1.277677108903695e+17, 1.277677108975571e+17, 1.27767710910682e+17, 1.27767710920682e+17, 1.277677109297445e+17, 1.277677109359945e+17, 1.27767710950682e+17, 1.27767710960682e+17, 1.27767710970682e+17, 1.27767710980682e+17, 1.27767710990682e+17, 1.27767711000682e+17, 1.277677110070883e+17, 1.277677110167757e+17, 1.27767711030682e+17, 1.27767711040682e+17, 1.27767711050682e+17, 1.27767711060682e+17, 1.277677110699008e+17, 1.27767711080682e+17, 1.27767711090682e+17, 1.27767711100682e+17, 1.27767711110682e+17, 1.277677111202132e+17, 1.27767711130682e+17, 1.27767711140682e+17, 1.27767711150682e+17, 1.27767711160682e+17, 1.27767711170057e+17, 1.27767711180682e+17, 1.27767711190682e+17, 1.27767711200682e+17, 1.27767711210682e+17, 1.277677112202132e+17, 1.27767711230682e+17, 1.27767711240682e+17, 1.27767711250682e+17, 1.27767711260682e+17, 1.277677112694319e+17, 1.27767711280682e+17, 1.27767711290682e+17, 1.27767711300682e+17, 1.27767711310682e+17, 1.277677113195882e+17, 1.27767711330682e+17, 1.27767711340682e+17, 1.27767711350682e+17, 1.27767711360682e+17, 1.27767711370682e+17, 1.277677113803695e+17, 1.27767711390682e+17, 1.27767711400682e+17, 1.27767711410682e+17, 1.27767711420682e+17, 1.277677114295882e+17, 1.27767711440682e+17, 1.27767711450682e+17, 1.27767711460682e+17, 1.27767711470682e+17, 1.277677114792756e+17, 1.27767711490682e+17, 1.27767711500682e+17, 1.27767711510682e+17, 1.27767711520682e+17, 1.277677115295882e+17, 1.27767711540682e+17, 1.27767711550682e+17, 1.27767711560682e+17, 1.27767711570682e+17, 1.277677115797445e+17, 1.27767711590682e+17, 1.27767711600682e+17, 1.27767711610682e+17, 1.27767711620682e+17, 1.277677116295884e+17, 1.27767711640682e+17, 1.27767711650682e+17, 1.27767711660682e+17, 1.27767711670682e+17, 1.277677116799008e+17, 1.27767711690682e+17, 1.27767711700682e+17, 1.27767711710682e+17, 1.27767711720682e+17, 1.27767711730057e+17, 1.277677117406821e+17, 1.27767711750682e+17, 1.27767711760682e+17, 1.27767711770682e+17, 1.277677117799007e+17, 1.27767711790682e+17, 1.27767711800682e+17, 1.27767711810682e+17, 1.27767711820682e+17, 1.277677118302132e+17, 1.27767711840682e+17, 1.27767711850682e+17, 1.27767711860682e+17, 1.27767711870682e+17, 1.277677118792758e+17, 1.27767711890682e+17, 1.27767711900682e+17, 1.27767711910682e+17, 1.27767711920682e+17, 1.27767711930682e+17, 1.27767711940682e+17, 1.27767711950682e+17, 1.27767711960682e+17, 1.27767711970682e+17, 1.277677119803695e+17, 1.277677119903695e+17, 1.277677120006821e+17, 1.27767712010682e+17, 1.27767712020682e+17, 1.27767712030682e+17, 1.277677120395884e+17, 1.27767712050682e+17, 1.27767712060682e+17, 1.27767712070682e+17, 1.27767712080682e+17, 1.277677120902132e+17, 1.27767712100682e+17, 1.27767712110682e+17, 1.27767712120682e+17, 1.27767712130682e+17, 1.277677121402132e+17, 1.27767712150682e+17, 1.27767712160682e+17, 1.27767712170682e+17, 1.27767712180682e+17, 1.277677121895882e+17, 1.27767712200682e+17, 1.27767712210682e+17, 1.27767712220682e+17, 1.27767712230682e+17, 1.277677122397445e+17, 1.27767712250682e+17, 1.27767712260682e+17, 1.27767712270682e+17, 1.27767712280682e+17, 1.277677122899008e+17, 1.27767712300682e+17, 1.27767712310682e+17, 1.27767712320682e+17, 1.27767712330682e+17, 1.277677123397445e+17, 1.27767712350682e+17, 1.27767712360682e+17, 1.277677123706821e+17, 1.27767712380682e+17, 1.27767712390057e+17, 1.27767712400682e+17, 1.27767712410682e+17, 1.27767712420682e+17, 1.27767712430682e+17, 1.277677124397444e+17, 1.27767712450682e+17, 1.27767712460682e+17, 1.27767712470682e+17, 1.277677124799007e+17, 1.27767712490682e+17, 1.27767712500682e+17, 1.27767712510682e+17, 1.27767712520057e+17, 1.27767712530682e+17, 1.27767712540682e+17, 1.27767712550682e+17, 1.27767712560057e+17, 1.27767712570682e+17, 1.27767712580682e+17, 1.27767712590682e+17, 1.277677126002132e+17, 1.27767712610682e+17, 1.27767712620682e+17, 1.277677126306821e+17, 1.277677126394319e+17, 1.27767712650682e+17, 1.27767712660682e+17, 1.27767712670682e+17, 1.277677126794319e+17, 1.27767712690682e+17, 1.27767712700682e+17, 1.27767712710682e+17, 1.277677127202132e+17, 1.27767712730682e+17, 1.27767712740682e+17, 1.27767712750682e+17, 1.277677127594321e+17, 1.27767712770682e+17, 1.27767712780682e+17, 1.27767712790682e+17, 1.277677127995884e+17, 1.27767712810682e+17, 1.27767712820682e+17, 1.27767712830682e+17, 1.277677128397445e+17, 1.27767712850682e+17, 1.27767712860682e+17, 1.27767712870682e+17, 1.277677128795882e+17, 1.277677128906821e+17, 1.27767712900682e+17, 1.27767712910682e+17, 1.277677129195882e+17, 1.27767712930682e+17, 1.27767712940682e+17, 1.27767712950682e+17, 1.277677129597444e+17, 1.27767712970682e+17, 1.27767712980682e+17, 1.27767712990682e+17, 1.277677129999007e+17, 1.27767713010682e+17, 1.27767713020682e+17, 1.27767713030682e+17, 1.277677130397445e+17, 1.27767713050682e+17, 1.27767713060682e+17, 1.27767713070682e+17, 1.277677130799008e+17, 1.27767713090682e+17, 1.27767713100682e+17, 1.27767713110682e+17, 1.277677131199008e+17, 1.27767713130682e+17, 1.27767713140682e+17, 1.27767713150682e+17, 1.27767713160057e+17, 1.27767713170682e+17, 1.27767713180682e+17, 1.27767713190682e+17, 1.277677131992758e+17, 1.27767713210682e+17, 1.27767713220682e+17, 1.27767713230682e+17, 1.277677132400571e+17, 1.27767713250682e+17, 1.277677132606821e+17, 1.27767713270682e+17, 1.277677132802132e+17, 1.27767713290682e+17, 1.27767713300682e+17, 1.27767713310682e+17, 1.277677133192758e+17, 1.27767713330682e+17, 1.27767713340682e+17, 1.27767713350682e+17, 1.277677133595882e+17, 1.27767713370682e+17, 1.27767713380682e+17, 1.27767713390682e+17, 1.277677133994319e+17, 1.27767713410682e+17, 1.27767713420682e+17, 1.27767713430682e+17, 1.277677134394321e+17, 1.27767713450682e+17, 1.27767713460682e+17, 1.27767713470682e+17, 1.277677134795882e+17, 1.27767713490682e+17, 1.27767713500682e+17, 1.27767713510682e+17, 1.277677135202132e+17, 1.27767713530682e+17, 1.27767713540682e+17, 1.27767713550682e+17, 1.277677135595884e+17, 1.27767713570682e+17, 1.27767713580682e+17, 1.27767713590682e+17, 1.277677135995882e+17, 1.27767713610682e+17, 1.27767713620682e+17, 1.27767713630682e+17, 1.277677136397445e+17, 1.27767713650682e+17, 1.27767713660682e+17, 1.27767713670682e+17, 1.277677136799008e+17, 1.27767713690682e+17, 1.27767713700682e+17, 1.27767713710682e+17, 1.277677137197445e+17, 1.27767713730682e+17, 1.27767713740682e+17, 1.27767713750682e+17, 1.277677137599007e+17, 1.27767713770682e+17, 1.277677137806821e+17, 1.27767713790682e+17, 1.27767713800057e+17, 1.27767713810682e+17, 1.27767713820682e+17, 1.27767713830682e+17, 1.277677138402132e+17, 1.27767713850682e+17, 1.27767713860682e+17, 1.27767713870682e+17, 1.27767713880057e+17, 1.27767713890682e+17, 1.27767713900682e+17, 1.27767713910682e+17, 1.277677139202132e+17, 1.27767713930682e+17, 1.27767713940682e+17, 1.27767713950682e+17, 1.277677139592758e+17, 1.27767713970682e+17, 1.27767713980682e+17, 1.27767713990682e+17, 1.277677139994321e+17, 1.27767714010682e+17, 1.27767714020682e+17, 1.27767714030682e+17, 1.277677140402132e+17, 1.27767714050682e+17, 1.27767714060682e+17, 1.27767714070682e+17, 1.277677140794319e+17, 1.27767714090682e+17, 1.27767714100682e+17, 1.27767714110682e+17, 1.27767714120057e+17, 1.27767714130682e+17, 1.27767714140682e+17, 1.27767714150682e+17, 1.277677141602132e+17, 1.27767714170682e+17, 1.27767714180682e+17, 1.27767714190682e+17, 1.277677141994319e+17, 1.27767714210682e+17, 1.27767714220682e+17, 1.27767714230682e+17, 1.277677142395882e+17, 1.27767714250682e+17, 1.27767714260682e+17, 1.27767714270682e+17, 1.277677142797445e+17, 1.27767714290682e+17, 1.27767714300682e+17, 1.27767714310682e+17, 1.277677143199008e+17, 1.27767714330682e+17, 1.27767714340682e+17, 1.27767714350682e+17, 1.277677143594319e+17, 1.27767714370682e+17, 1.27767714380682e+17, 1.27767714390682e+17, 1.277677143997445e+17, 1.277677144106821e+17, 1.27767714420682e+17, 1.27767714430682e+17, 1.277677144399008e+17, 1.27767714450682e+17, 1.27767714460682e+17, 1.27767714470682e+17, 1.277677144800571e+17, 1.27767714490682e+17, 1.27767714500682e+17, 1.27767714510682e+17, 1.277677145194321e+17, 1.27767714530682e+17, 1.27767714540682e+17, 1.27767714550682e+17, 1.27767714560057e+17, 1.27767714570682e+17, 1.27767714580682e+17, 1.27767714590682e+17, 1.277677146002132e+17, 1.27767714610682e+17, 1.27767714620682e+17, 1.27767714630682e+17, 1.277677146392758e+17, 1.27767714650682e+17, 1.27767714660682e+17, 1.277677146706821e+17, 1.277677146794319e+17, 1.27767714690682e+17, 1.27767714700682e+17, 1.27767714710682e+17, 1.277677147202132e+17, 1.27767714730682e+17, 1.27767714740682e+17, 1.27767714750682e+17, 1.277677147592758e+17, 1.27767714770682e+17, 1.27767714780682e+17, 1.27767714790682e+17, 1.277677147994321e+17, 1.27767714810682e+17, 1.27767714820682e+17, 1.27767714830682e+17, 1.277677148395884e+17, 1.27767714850682e+17, 1.27767714860682e+17, 1.27767714870682e+17, 1.277677148794319e+17, 1.27767714890682e+17, 1.27767714900682e+17, 1.27767714910682e+17, 1.277677149195882e+17, 1.277677149306821e+17, 1.27767714940682e+17, 1.277677149486508e+17, 1.277677149586508e+17, 1.27767714970682e+17, 1.27767714980682e+17, 1.27767714990682e+17, 1.277677149999008e+17, 1.27767715010682e+17, 1.27767715020682e+17, 1.27767715030682e+17, 1.277677150395884e+17, 1.27767715050682e+17, 1.27767715060682e+17, 1.27767715070682e+17, 1.277677150797445e+17, 1.27767715090682e+17, 1.27767715100682e+17, 1.27767715110682e+17, 1.277677151199008e+17, 1.27767715130682e+17, 1.27767715140682e+17, 1.27767715150682e+17, 1.27767715160057e+17, 1.27767715170682e+17, 1.27767715180682e+17, 1.27767715190682e+17, 1.277677151999008e+17, 1.27767715210682e+17, 1.27767715220682e+17, 1.27767715230682e+17, 1.277677152399008e+17, 1.27767715250682e+17, 1.27767715260682e+17, 1.27767715270682e+17, 1.277677152799007e+17, 1.27767715290682e+17, 1.277677153006821e+17, 1.27767715310682e+17, 1.27767715320057e+17, 1.27767715330682e+17, 1.27767715340682e+17, 1.27767715350682e+17, 1.277677153602132e+17, 1.27767715370682e+17, 1.27767715380682e+17, 1.27767715390682e+17, 1.277677153992758e+17, 1.27767715410682e+17, 1.27767715420682e+17, 1.27767715430682e+17, 1.277677154394319e+17, 1.27767715450682e+17, 1.27767715460682e+17, 1.27767715470682e+17, 1.277677154800571e+17, 1.27767715490682e+17, 1.27767715500682e+17, 1.27767715510682e+17, 1.277677155194321e+17, 1.27767715530682e+17, 1.27767715540682e+17, 1.27767715550682e+17, 1.277677155595884e+17, 1.27767715570682e+17, 1.27767715580682e+17, 1.27767715590682e+17, 1.277677155997445e+17, 1.27767715610682e+17, 1.27767715620682e+17, 1.27767715630682e+17, 1.277677156397445e+17, 1.27767715650682e+17, 1.27767715660682e+17, 1.27767715670682e+17, 1.277677156795882e+17, 1.27767715690682e+17, 1.27767715700682e+17, 1.27767715710682e+17, 1.277677157197445e+17, 1.27767715730682e+17, 1.27767715740682e+17, 1.27767715750682e+17, 1.277677157599008e+17, 1.27767715770682e+17, 1.27767715780682e+17, 1.27767715790682e+17, 1.27767715800682e+17, 1.27767715810682e+17, 1.277677158206821e+17, 1.27767715830682e+17, 1.277677158399008e+17, 1.27767715850682e+17, 1.27767715860682e+17, 1.27767715870682e+17, 1.27767715880057e+17, 1.27767715890682e+17, 1.27767715900682e+17, 1.27767715910682e+17, 1.277677159202132e+17, 1.27767715930682e+17, 1.27767715940682e+17, 1.27767715950682e+17, 1.277677159597445e+17, 1.27767715970682e+17, 1.27767715980682e+17, 1.27767715990682e+17, 1.277677160000571e+17, 1.27767716010682e+17, 1.27767716020682e+17, 1.27767716030682e+17, 1.277677160402132e+17, 1.27767716050682e+17, 1.27767716060682e+17, 1.27767716070682e+17, 1.277677160794321e+17, 1.27767716090682e+17, 1.27767716100682e+17, 1.27767716110682e+17, 1.277677161195884e+17, 1.27767716130682e+17, 1.27767716140682e+17, 1.27767716150682e+17, 1.277677161592758e+17, 1.27767716170682e+17, 1.27767716180682e+17, 1.277677161906821e+17, 1.277677161994319e+17, 1.27767716210682e+17, 1.27767716220682e+17, 1.27767716230682e+17, 1.277677162395882e+17, 1.27767716250682e+17, 1.27767716260682e+17, 1.27767716270682e+17, 1.277677162797445e+17, 1.27767716290682e+17, 1.27767716300682e+17, 1.27767716310682e+17, 1.277677163203695e+17, 1.27767716330682e+17, 1.27767716340682e+17, 1.27767716350682e+17, 1.277677163595882e+17, 1.27767716370682e+17, 1.27767716380682e+17, 1.27767716390682e+17, 1.277677164005257e+17, 1.27767716410682e+17, 1.27767716420682e+17, 1.27767716430682e+17, 1.277677164399008e+17, 1.277677164506821e+17, 1.27767716460682e+17, 1.27767716470682e+17, 1.277677164799008e+17, 1.27767716490682e+17, 1.27767716500682e+17, 1.27767716510682e+17, 1.277677165200571e+17, 1.27767716530682e+17, 1.27767716540682e+17, 1.27767716550682e+17, 1.277677165597445e+17, 1.27767716570682e+17, 1.27767716580682e+17, 1.27767716590682e+17, 1.27767716600057e+17, 1.27767716610682e+17, 1.27767716620682e+17, 1.27767716630682e+17, 1.277677166402132e+17, 1.27767716650682e+17, 1.27767716660682e+17, 1.27767716670682e+17, 1.277677166792758e+17, 1.27767716690682e+17, 1.27767716700682e+17, 1.277677167106821e+17, 1.277677167194319e+17, 1.27767716730682e+17, 1.27767716740682e+17, 1.27767716750682e+17, 1.277677167602132e+17, 1.27767716770682e+17, 1.27767716780682e+17, 1.27767716790682e+17, 1.277677167992758e+17, 1.27767716810682e+17, 1.27767716820682e+17, 1.27767716830682e+17, 1.277677168394321e+17, 1.27767716850682e+17, 1.27767716860682e+17, 1.27767716870682e+17, 1.277677168795884e+17, 1.27767716890682e+17, 1.27767716900682e+17, 1.27767716910682e+17, 1.277677169202132e+17, 1.27767716930682e+17, 1.27767716940682e+17, 1.27767716950682e+17, 1.277677169594319e+17, 1.27767716970682e+17, 1.27767716980682e+17, 1.27767716990682e+17, 1.277677169995882e+17, 1.27767717010682e+17, 1.27767717020682e+17, 1.27767717030682e+17, 1.277677170397444e+17, 1.27767717050682e+17, 1.27767717060682e+17, 1.27767717070682e+17, 1.277677170794321e+17, 1.27767717090682e+17, 1.27767717100682e+17, 1.27767717110682e+17, 1.277677171197445e+17, 1.27767717130682e+17, 1.27767717140682e+17, 1.27767717150682e+17, 1.277677171599008e+17, 1.27767717170682e+17, 1.27767717180682e+17, 1.27767717190682e+17, 1.27767717200057e+17, 1.27767717210682e+17, 1.27767717220682e+17, 1.27767717230682e+17, 1.27767717240057e+17, 1.27767717250682e+17, 1.27767717260682e+17, 1.27767717270682e+17, 1.277677172797445e+17, 1.27767717290682e+17, 1.27767717300682e+17, 1.27767717310682e+17, 1.277677173200571e+17, 1.27767717330682e+17, 1.277677173406821e+17, 1.27767717350682e+17, 1.277677173602132e+17, 1.27767717370682e+17, 1.27767717380682e+17, 1.27767717390682e+17, 1.277677173992758e+17, 1.27767717410682e+17, 1.27767717420682e+17, 1.27767717430682e+17, 1.27767717440057e+17, 1.27767717450682e+17, 1.27767717460682e+17, 1.27767717470682e+17, 1.277677174802131e+17, 1.27767717490682e+17, 1.27767717500682e+17, 1.27767717510682e+17, 1.277677175194321e+17, 1.27767717530682e+17, 1.27767717540682e+17, 1.27767717550682e+17, 1.277677175602132e+17, 1.27767717570682e+17, 1.27767717580682e+17, 1.27767717590682e+17, 1.277677176002132e+17, 1.27767717610682e+17, 1.27767717620682e+17, 1.27767717630682e+17, 1.277677176392756e+17, 1.27767717650682e+17, 1.27767717660682e+17, 1.27767717670682e+17, 1.277677176795882e+17, 1.27767717690682e+17, 1.27767717700682e+17, 1.27767717710682e+17, 1.277677177197445e+17, 1.27767717730682e+17, 1.27767717740682e+17, 1.27767717750682e+17, 1.277677177599008e+17, 1.27767717770682e+17, 1.27767717780682e+17, 1.27767717790682e+17, 1.277677177999008e+17, 1.27767717810682e+17, 1.27767717820682e+17, 1.27767717830682e+17, 1.277677178397445e+17, 1.27767717850682e+17, 1.27767717860682e+17, 1.27767717870682e+17, 1.277677178799008e+17, 1.27767717890682e+17, 1.27767717900682e+17, 1.27767717910682e+17, 1.27767717920057e+17, 1.27767717930682e+17, 1.27767717940682e+17, 1.27767717950682e+17, 1.27767717960682e+17, 1.27767717970682e+17, 1.27767717980682e+17, 1.27767717990682e+17, 1.27767718000682e+17, 1.27767718010682e+17, 1.27767718020682e+17, 1.27767718030682e+17, 1.277677180391195e+17, 1.277677180480257e+17, 1.27767718060682e+17, 1.27767718070682e+17, 1.27767718080682e+17, 1.27767718090682e+17, 1.27767718100682e+17, 1.277677181092758e+17, 1.277677181183383e+17, 1.27767718130682e+17, 1.27767718140682e+17, 1.277677181494321e+17, 1.27767718160682e+17, 1.27767718168182e+17, 1.27767718180682e+17, 1.277677181872445e+17, 1.27767718200682e+17, 1.27767718210682e+17, 1.277677182192758e+17, 1.277677182306821e+17, 1.277677182374008e+17, 1.277677182464634e+17, 1.27767718260682e+17, 1.27767718270682e+17, 1.277677182794319e+17, 1.27767718290682e+17, 1.277677182974007e+17, 1.277677183066195e+17, 1.27767718320682e+17, 1.27767718330682e+17, 1.277677183394321e+17},
			             {1.27767684410682e+17, 1.27767684420682e+17, 1.27767684430682e+17, 1.27767684440682e+17, 1.27767684450682e+17, 1.27767684460682e+17, 1.27767684470682e+17, 1.277676844806821e+17, 1.27767684490682e+17, 1.27767684500682e+17, 1.27767684510682e+17, 1.27767684520682e+17, 1.27767684530682e+17, 1.27767684540682e+17, 1.27767684550682e+17, 1.27767684560682e+17, 1.27767684570682e+17, 1.27767684580682e+17, 1.27767684590682e+17, 1.27767684600682e+17, 1.27767684610682e+17, 1.27767684620682e+17, 1.27767684630682e+17, 1.27767684640682e+17, 1.27767684650682e+17, 1.27767684660682e+17, 1.27767684670682e+17, 1.27767684680682e+17, 1.27767684690682e+17, 1.27767684700682e+17, 1.27767684710682e+17, 1.27767684720682e+17, 1.27767684730682e+17, 1.277676847406821e+17, 1.27767684750682e+17, 1.27767684760682e+17, 1.27767684770682e+17, 1.27767684780682e+17, 1.27767684790682e+17, 1.27767684800682e+17, 1.27767684810682e+17, 1.27767684820682e+17, 1.27767684830682e+17, 1.27767684840682e+17, 1.27767684850682e+17, 1.27767684860682e+17, 1.27767684870682e+17, 1.27767684880682e+17, 1.27767684890682e+17, 1.27767684900682e+17, 1.27767684910682e+17, 1.27767684920682e+17, 1.27767684930682e+17, 1.27767684940682e+17, 1.27767684950682e+17, 1.27767684960682e+17, 1.27767684970682e+17, 1.27767684980682e+17, 1.27767684990682e+17, 1.277676850006821e+17, 1.27767685010682e+17, 1.27767685020682e+17, 1.27767685030682e+17, 1.27767685040682e+17, 1.27767685050682e+17, 1.27767685060682e+17, 1.27767685070682e+17, 1.27767685080682e+17, 1.27767685090682e+17, 1.27767685100682e+17, 1.27767685110682e+17, 1.27767685120682e+17, 1.27767685130682e+17, 1.27767685140682e+17, 1.27767685150682e+17, 1.27767685160682e+17, 1.27767685170682e+17, 1.27767685180682e+17, 1.27767685190682e+17, 1.27767685200682e+17, 1.27767685210682e+17, 1.27767685220682e+17, 1.27767685230682e+17, 1.27767685240682e+17, 1.27767685250682e+17, 1.27767685260682e+17, 1.27767685270682e+17, 1.27767685280682e+17, 1.27767685290682e+17, 1.27767685300682e+17, 1.27767685310682e+17, 1.27767685320682e+17, 1.27767685330682e+17, 1.27767685340682e+17, 1.27767685350682e+17, 1.27767685360682e+17, 1.277676853706821e+17, 1.27767685380682e+17, 1.27767685390682e+17, 1.27767685400682e+17, 1.27767685410682e+17, 1.27767685420682e+17, 1.27767685430682e+17, 1.27767685440682e+17, 1.27767685450682e+17, 1.27767685460682e+17, 1.27767685470682e+17, 1.27767685480682e+17, 1.27767685490682e+17, 1.27767685500682e+17, 1.27767685510682e+17, 1.27767685520682e+17, 1.27767685530682e+17, 1.27767685540682e+17, 1.27767685550682e+17, 1.27767685560682e+17, 1.27767685570682e+17, 1.27767685580682e+17, 1.27767685590682e+17, 1.27767685600682e+17, 1.27767685610682e+17, 1.27767685620682e+17, 1.277676856306821e+17, 1.27767685640682e+17, 1.27767685650682e+17, 1.27767685660682e+17, 1.27767685670682e+17, 1.27767685680682e+17, 1.27767685690682e+17, 1.27767685700682e+17, 1.27767685710682e+17, 1.27767685720682e+17, 1.27767685730682e+17, 1.27767685740682e+17, 1.27767685750682e+17, 1.27767685760682e+17, 1.27767685770682e+17, 1.27767685780682e+17, 1.27767685790682e+17, 1.27767685800682e+17, 1.27767685810682e+17, 1.27767685820682e+17, 1.27767685830682e+17, 1.27767685840682e+17, 1.27767685850682e+17, 1.27767685860682e+17, 1.27767685870682e+17, 1.27767685880682e+17, 1.277676858906821e+17, 1.27767685900682e+17, 1.27767685910682e+17, 1.27767685920682e+17, 1.27767685930682e+17, 1.27767685940682e+17, 1.27767685950682e+17, 1.27767685960682e+17, 1.27767685970682e+17, 1.27767685980682e+17, 1.27767685990682e+17, 1.27767686000682e+17, 1.27767686010682e+17, 1.27767686020682e+17, 1.27767686030682e+17, 1.27767686040682e+17, 1.27767686050682e+17, 1.27767686060682e+17, 1.27767686070682e+17, 1.27767686080682e+17, 1.27767686090682e+17, 1.27767686100682e+17, 1.27767686110682e+17, 1.27767686120682e+17, 1.27767686130682e+17, 1.27767686140682e+17, 1.27767686150682e+17, 1.27767686160682e+17, 1.27767686170682e+17, 1.27767686180682e+17, 1.27767686190682e+17, 1.27767686200682e+17, 1.27767686210682e+17, 1.27767686220682e+17, 1.27767686230682e+17, 1.27767686240682e+17, 1.27767686250682e+17, 1.277676862606821e+17, 1.27767686270682e+17, 1.27767686280682e+17, 1.27767686290682e+17, 1.27767686300682e+17, 1.27767686310682e+17, 1.27767686320682e+17, 1.27767686330682e+17, 1.27767686340682e+17, 1.27767686350682e+17, 1.27767686360682e+17, 1.27767686370682e+17, 1.27767686380682e+17, 1.27767686390682e+17, 1.27767686400682e+17, 1.27767686410682e+17, 1.27767686420682e+17, 1.27767686430682e+17, 1.27767686440682e+17, 1.27767686450682e+17, 1.27767686460682e+17, 1.27767686470682e+17, 1.27767686480682e+17, 1.27767686490682e+17, 1.27767686500682e+17, 1.27767686510682e+17, 1.277676865206821e+17, 1.27767686530682e+17, 1.27767686540682e+17, 1.27767686550682e+17, 1.27767686560682e+17, 1.27767686570682e+17, 1.27767686580682e+17, 1.27767686590682e+17, 1.27767686600682e+17, 1.27767686610682e+17, 1.27767686620682e+17, 1.27767686630682e+17, 1.27767686640682e+17, 1.27767686650682e+17, 1.27767686660682e+17, 1.27767686670682e+17, 1.27767686680682e+17, 1.27767686690682e+17, 1.27767686700682e+17, 1.27767686710682e+17, 1.27767686720682e+17, 1.27767686730682e+17, 1.27767686740682e+17, 1.27767686750682e+17, 1.27767686760682e+17, 1.27767686770682e+17, 1.277676867806821e+17, 1.27767686790682e+17, 1.27767686800682e+17, 1.27767686810682e+17, 1.27767686820682e+17, 1.27767686830682e+17, 1.27767686840682e+17, 1.27767686850682e+17, 1.27767686860682e+17, 1.27767686870682e+17, 1.27767686880682e+17, 1.27767686890682e+17, 1.27767686900682e+17, 1.27767686910682e+17, 1.27767686920682e+17, 1.27767686930682e+17, 1.27767686940682e+17, 1.27767686950682e+17, 1.27767686960682e+17, 1.27767686970682e+17, 1.27767686980682e+17, 1.27767686990682e+17, 1.27767687000682e+17, 1.27767687010682e+17, 1.27767687020682e+17, 1.27767687030682e+17, 1.27767687040682e+17, 1.27767687050682e+17, 1.27767687060682e+17, 1.27767687070682e+17, 1.27767687080682e+17, 1.27767687090682e+17, 1.27767687100682e+17, 1.27767687110682e+17},
			             {1.27767694480682e+17, 1.27767694490682e+17, 1.27767694500682e+17, 1.27767694510682e+17, 1.27767694520682e+17, 1.27767694530682e+17, 1.27767694540682e+17, 1.27767694550682e+17, 1.27767694560682e+17, 1.27767694570682e+17, 1.27767694580682e+17, 1.27767694590682e+17, 1.27767694600682e+17, 1.27767694610682e+17, 1.27767694620682e+17, 1.27767694630682e+17, 1.27767694640682e+17, 1.27767694650682e+17, 1.27767694660682e+17, 1.27767694670682e+17, 1.277676946806821e+17, 1.27767694690682e+17, 1.27767694700682e+17, 1.27767694710682e+17, 1.27767694720682e+17, 1.27767694730682e+17, 1.27767694740682e+17, 1.27767694750682e+17, 1.27767694760682e+17, 1.27767694770682e+17, 1.27767694780682e+17, 1.27767694790682e+17, 1.27767694800682e+17, 1.27767694810682e+17, 1.27767694820682e+17, 1.27767694830682e+17, 1.27767694840682e+17, 1.27767694850682e+17, 1.27767694860682e+17, 1.27767694870682e+17, 1.27767694880682e+17, 1.27767694890682e+17, 1.27767694900682e+17, 1.27767694910682e+17, 1.27767694920682e+17, 1.27767694930682e+17, 1.27767694940682e+17, 1.27767694950682e+17, 1.27767694960682e+17, 1.27767694970682e+17, 1.27767694980682e+17, 1.27767694990682e+17, 1.27767695000682e+17, 1.27767695010682e+17, 1.27767695020682e+17, 1.27767695030682e+17, 1.27767695040682e+17, 1.277676950506821e+17, 1.27767695060682e+17, 1.27767695070682e+17, 1.27767695080682e+17, 1.27767695090682e+17, 1.27767695100682e+17, 1.27767695110682e+17, 1.27767695120682e+17, 1.27767695130682e+17, 1.27767695140682e+17, 1.27767695150682e+17, 1.27767695160682e+17, 1.27767695170682e+17, 1.27767695180682e+17, 1.27767695190682e+17, 1.27767695200682e+17, 1.27767695210682e+17, 1.27767695220682e+17, 1.27767695230682e+17, 1.27767695240682e+17, 1.27767695250682e+17, 1.27767695260682e+17, 1.27767695270682e+17, 1.27767695280682e+17, 1.27767695290682e+17, 1.27767695300682e+17, 1.277676953106821e+17, 1.27767695320682e+17, 1.27767695330682e+17, 1.27767695340682e+17, 1.27767695350682e+17, 1.27767695360682e+17, 1.27767695370682e+17, 1.27767695380682e+17, 1.27767695390682e+17, 1.27767695400682e+17, 1.27767695410682e+17, 1.27767695420682e+17, 1.27767695430682e+17, 1.27767695440682e+17, 1.27767695450682e+17, 1.27767695460682e+17, 1.27767695470682e+17, 1.27767695480682e+17, 1.27767695490682e+17, 1.27767695500682e+17, 1.27767695510682e+17, 1.27767695520682e+17, 1.27767695530682e+17, 1.27767695540682e+17, 1.27767695550682e+17, 1.27767695560682e+17, 1.277676955706821e+17, 1.27767695580682e+17, 1.27767695590682e+17, 1.27767695600682e+17, 1.27767695610682e+17, 1.27767695620682e+17, 1.27767695630682e+17, 1.27767695640682e+17, 1.27767695650682e+17, 1.27767695660682e+17, 1.27767695670682e+17, 1.27767695680682e+17, 1.27767695690682e+17, 1.27767695700682e+17, 1.27767695710682e+17, 1.27767695720682e+17, 1.27767695730682e+17, 1.27767695740682e+17, 1.27767695750682e+17, 1.27767695760682e+17, 1.27767695770682e+17, 1.27767695780682e+17, 1.27767695790682e+17, 1.27767695800682e+17, 1.27767695810682e+17, 1.27767695820682e+17, 1.27767695830682e+17, 1.27767695840682e+17, 1.27767695850682e+17, 1.27767695860682e+17, 1.27767695870682e+17, 1.27767695880682e+17, 1.27767695890682e+17, 1.27767695900682e+17, 1.27767695910682e+17, 1.27767695920682e+17, 1.27767695930682e+17, 1.277676959406821e+17, 1.27767695950682e+17, 1.27767695960682e+17, 1.27767695970682e+17, 1.27767695980682e+17, 1.27767695990682e+17, 1.27767696000682e+17, 1.27767696010682e+17, 1.27767696020682e+17, 1.27767696030682e+17, 1.27767696040682e+17, 1.27767696050682e+17, 1.27767696060682e+17, 1.27767696070682e+17, 1.27767696080682e+17, 1.27767696090682e+17, 1.27767696100682e+17, 1.27767696110682e+17, 1.27767696120682e+17, 1.27767696130682e+17, 1.27767696140682e+17, 1.27767696150682e+17, 1.27767696160682e+17, 1.27767696170682e+17, 1.27767696180682e+17, 1.27767696190682e+17, 1.277676962006821e+17, 1.27767696210682e+17, 1.27767696220682e+17, 1.27767696230682e+17, 1.27767696240682e+17, 1.27767696250682e+17, 1.27767696260682e+17, 1.27767696270682e+17, 1.27767696280682e+17, 1.27767696290682e+17, 1.27767696300682e+17, 1.27767696310682e+17, 1.27767696320682e+17, 1.27767696330682e+17, 1.27767696340682e+17, 1.27767696350682e+17, 1.27767696360682e+17, 1.27767696370682e+17, 1.27767696380682e+17, 1.27767696390682e+17, 1.27767696400682e+17, 1.27767696410682e+17, 1.27767696420682e+17, 1.27767696430682e+17, 1.27767696440682e+17, 1.27767696450682e+17, 1.277676964606821e+17, 1.27767696470682e+17, 1.27767696480682e+17, 1.27767696490682e+17, 1.27767696500682e+17, 1.27767696510682e+17, 1.27767696520682e+17, 1.27767696530682e+17, 1.27767696540682e+17, 1.27767696550682e+17, 1.27767696560682e+17, 1.27767696570682e+17, 1.27767696580682e+17, 1.27767696590682e+17, 1.27767696600682e+17, 1.27767696610682e+17, 1.27767696620682e+17, 1.27767696630682e+17, 1.27767696640682e+17, 1.27767696650682e+17, 1.27767696660682e+17, 1.27767696670682e+17, 1.27767696680682e+17, 1.27767696690682e+17, 1.27767696700682e+17, 1.27767696710682e+17, 1.27767696720682e+17, 1.27767696730682e+17, 1.27767696740682e+17, 1.27767696750682e+17, 1.27767696760682e+17, 1.27767696770682e+17, 1.27767696780682e+17, 1.27767696790682e+17, 1.27767696800682e+17, 1.27767696810682e+17, 1.27767696820682e+17, 1.277676968306821e+17, 1.27767696840682e+17, 1.27767696850682e+17, 1.27767696860682e+17, 1.27767696870682e+17, 1.27767696880682e+17, 1.27767696890682e+17, 1.27767696900682e+17, 1.27767696910682e+17, 1.27767696920682e+17, 1.27767696930682e+17, 1.27767696940682e+17, 1.27767696950682e+17, 1.27767696960682e+17, 1.27767696970682e+17, 1.27767696980682e+17, 1.27767696990682e+17, 1.27767697000682e+17, 1.27767697010682e+17, 1.27767697020682e+17, 1.27767697030682e+17, 1.27767697040682e+17, 1.27767697050682e+17, 1.27767697060682e+17, 1.27767697070682e+17, 1.27767697080682e+17, 1.277676970906821e+17, 1.27767697100682e+17, 1.27767697110682e+17, 1.27767697120682e+17, 1.27767697130682e+17, 1.27767697140682e+17, 1.27767697150682e+17, 1.27767697160682e+17, 1.27767697170682e+17, 1.27767697180682e+17, 1.27767697190682e+17, 1.27767697200682e+17, 1.27767697210682e+17, 1.27767697220682e+17, 1.27767697230682e+17, 1.27767697240682e+17, 1.27767697250682e+17, 1.27767697260682e+17, 1.27767697270682e+17, 1.27767697280682e+17, 1.27767697290682e+17, 1.27767697300682e+17, 1.27767697310682e+17, 1.27767697320682e+17, 1.27767697330682e+17, 1.27767697340682e+17, 1.277676973506821e+17, 1.27767697360682e+17, 1.27767697370682e+17, 1.27767697380682e+17, 1.27767697390682e+17, 1.27767697400682e+17, 1.27767697410682e+17, 1.27767697420682e+17, 1.27767697430682e+17, 1.27767697440682e+17, 1.27767697450682e+17, 1.27767697460682e+17, 1.27767697470682e+17, 1.27767697480682e+17, 1.27767697490682e+17, 1.27767697500682e+17, 1.27767697510682e+17, 1.27767697520682e+17, 1.27767697530682e+17, 1.27767697540682e+17, 1.27767697550682e+17, 1.27767697560682e+17, 1.27767697570682e+17, 1.27767697580682e+17, 1.27767697590682e+17, 1.27767697600682e+17, 1.27767697610682e+17, 1.27767697620682e+17, 1.27767697630682e+17, 1.27767697640682e+17, 1.27767697650682e+17, 1.27767697660682e+17, 1.27767697670682e+17, 1.27767697680682e+17, 1.27767697690682e+17, 1.27767697700682e+17, 1.27767697710682e+17, 1.27767697720682e+17, 1.27767697730682e+17, 1.27767697740682e+17, 1.27767697750682e+17, 1.27767697760682e+17, 1.27767697770682e+17, 1.27767697780682e+17, 1.27767697790682e+17, 1.27767697800682e+17, 1.27767697810682e+17, 1.27767697820682e+17, 1.27767697830682e+17, 1.27767697840682e+17, 1.27767697850682e+17, 1.27767697860682e+17, 1.27767697870682e+17, 1.27767697880682e+17, 1.27767697890682e+17, 1.27767697900682e+17, 1.27767697910682e+17, 1.27767697920682e+17, 1.27767697930682e+17, 1.27767697940682e+17, 1.27767697950682e+17, 1.27767697960682e+17, 1.27767697970682e+17, 1.277676979806821e+17, 1.27767697990682e+17, 1.27767698000682e+17, 1.27767698010682e+17, 1.27767698020682e+17, 1.27767698030682e+17, 1.27767698040682e+17, 1.27767698050682e+17, 1.27767698060682e+17, 1.27767698070682e+17, 1.27767698080682e+17, 1.27767698090682e+17, 1.27767698100682e+17, 1.27767698110682e+17, 1.27767698120682e+17, 1.27767698130682e+17, 1.27767698140682e+17, 1.27767698150682e+17, 1.27767698160682e+17, 1.27767698170682e+17, 1.27767698180682e+17, 1.27767698190682e+17, 1.27767698200682e+17, 1.27767698210682e+17, 1.27767698220682e+17, 1.27767698230682e+17, 1.277676982406821e+17, 1.27767698250682e+17, 1.27767698260682e+17, 1.27767698270682e+17, 1.27767698280682e+17, 1.27767698290682e+17, 1.27767698300682e+17, 1.27767698310682e+17, 1.27767698320682e+17, 1.27767698330682e+17, 1.27767698340682e+17, 1.27767698350682e+17, 1.27767698360682e+17, 1.27767698370682e+17, 1.27767698380682e+17, 1.27767698390682e+17, 1.27767698400682e+17, 1.27767698410682e+17, 1.27767698420682e+17, 1.27767698430682e+17, 1.27767698440682e+17, 1.27767698450682e+17, 1.27767698460682e+17, 1.27767698470682e+17, 1.27767698480682e+17, 1.27767698490682e+17, 1.277676985006821e+17, 1.27767698510682e+17, 1.27767698520682e+17, 1.27767698530682e+17, 1.27767698540682e+17, 1.27767698550682e+17, 1.27767698560682e+17, 1.27767698570682e+17, 1.27767698580682e+17, 1.27767698590682e+17, 1.27767698600682e+17, 1.27767698610682e+17, 1.27767698620682e+17, 1.27767698630682e+17, 1.27767698640682e+17, 1.27767698650682e+17, 1.27767698660682e+17, 1.27767698670682e+17, 1.27767698680682e+17, 1.27767698690682e+17, 1.27767698700682e+17, 1.27767698710682e+17, 1.27767698720682e+17, 1.27767698730682e+17, 1.27767698740682e+17, 1.27767698750682e+17, 1.27767698760682e+17, 1.27767698770682e+17, 1.27767698780682e+17, 1.27767698790682e+17, 1.27767698800682e+17, 1.27767698810682e+17, 1.27767698820682e+17, 1.27767698830682e+17, 1.27767698840682e+17, 1.27767698850682e+17, 1.27767698860682e+17, 1.277676988706821e+17, 1.27767698880682e+17, 1.27767698890682e+17, 1.27767698900682e+17, 1.27767698910682e+17, 1.27767698920682e+17, 1.27767698930682e+17, 1.27767698940682e+17, 1.27767698950682e+17, 1.27767698960682e+17, 1.27767698970682e+17, 1.27767698980682e+17, 1.27767698990682e+17, 1.27767699000682e+17, 1.27767699010682e+17, 1.27767699020682e+17, 1.27767699030682e+17, 1.27767699040682e+17, 1.27767699050682e+17, 1.27767699060682e+17, 1.27767699070682e+17, 1.27767699080682e+17},
			             {1.27767691460682e+17, 1.27767691470682e+17, 1.27767691480682e+17, 1.277676914906821e+17, 1.27767691500682e+17, 1.27767691510682e+17, 1.27767691520682e+17, 1.27767691530682e+17, 1.27767691540682e+17, 1.27767691550682e+17, 1.27767691560682e+17, 1.27767691570682e+17, 1.27767691580682e+17, 1.27767691590682e+17, 1.27767691600682e+17, 1.27767691610682e+17, 1.27767691620682e+17, 1.27767691630682e+17, 1.27767691640682e+17, 1.27767691650682e+17, 1.27767691660682e+17, 1.27767691670682e+17, 1.27767691680682e+17, 1.27767691690682e+17, 1.27767691700682e+17, 1.27767691710682e+17, 1.27767691720682e+17, 1.27767691730682e+17, 1.27767691740682e+17, 1.277676917506821e+17, 1.27767691760682e+17, 1.27767691770682e+17, 1.27767691780682e+17, 1.27767691790682e+17, 1.27767691800682e+17, 1.27767691810682e+17, 1.27767691820682e+17, 1.27767691830682e+17, 1.27767691840682e+17, 1.27767691850682e+17, 1.27767691860682e+17, 1.27767691870682e+17, 1.27767691880682e+17, 1.27767691890682e+17, 1.27767691900682e+17, 1.27767691910682e+17, 1.27767691920682e+17, 1.27767691930682e+17, 1.27767691940682e+17, 1.27767691950682e+17, 1.27767691960682e+17, 1.27767691970682e+17, 1.27767691980682e+17, 1.27767691990682e+17, 1.27767692000682e+17, 1.27767692010682e+17, 1.27767692020682e+17, 1.27767692030682e+17, 1.27767692040682e+17, 1.27767692050682e+17, 1.27767692060682e+17, 1.27767692070682e+17, 1.27767692080682e+17, 1.27767692090682e+17, 1.27767692100682e+17, 1.27767692110682e+17, 1.277676921206821e+17, 1.27767692130682e+17, 1.27767692140682e+17, 1.27767692150682e+17, 1.27767692160682e+17, 1.27767692170682e+17, 1.27767692180682e+17, 1.27767692190682e+17, 1.27767692200682e+17, 1.27767692210682e+17, 1.27767692220682e+17, 1.27767692230682e+17, 1.27767692240682e+17, 1.27767692250682e+17, 1.27767692260682e+17, 1.27767692270682e+17, 1.27767692280682e+17, 1.27767692290682e+17, 1.27767692300682e+17, 1.27767692310682e+17, 1.27767692320682e+17, 1.27767692330682e+17, 1.27767692340682e+17, 1.27767692350682e+17, 1.27767692360682e+17, 1.27767692370682e+17, 1.277676923806821e+17, 1.27767692390682e+17, 1.27767692400682e+17, 1.27767692410682e+17, 1.27767692420682e+17, 1.27767692430682e+17, 1.27767692440682e+17, 1.27767692450682e+17, 1.27767692460682e+17, 1.27767692470682e+17, 1.27767692480682e+17, 1.27767692490682e+17, 1.27767692500682e+17, 1.27767692510682e+17, 1.27767692520682e+17, 1.27767692530682e+17, 1.27767692540682e+17, 1.27767692550682e+17, 1.27767692560682e+17, 1.27767692570682e+17, 1.27767692580682e+17, 1.27767692590682e+17, 1.27767692600682e+17, 1.27767692610682e+17, 1.27767692620682e+17, 1.27767692630682e+17, 1.277676926406821e+17, 1.27767692650682e+17, 1.27767692660682e+17, 1.27767692670682e+17, 1.27767692680682e+17, 1.27767692690682e+17, 1.27767692700682e+17, 1.27767692710682e+17, 1.27767692720682e+17, 1.27767692730682e+17, 1.27767692740682e+17, 1.27767692750682e+17, 1.27767692760682e+17, 1.27767692770682e+17, 1.27767692780682e+17, 1.27767692790682e+17, 1.27767692800682e+17, 1.27767692810682e+17, 1.27767692820682e+17, 1.27767692830682e+17, 1.27767692840682e+17, 1.27767692850682e+17, 1.27767692860682e+17, 1.27767692870682e+17, 1.27767692880682e+17, 1.27767692890682e+17, 1.27767692900682e+17, 1.27767692910682e+17, 1.27767692920682e+17, 1.27767692930682e+17, 1.27767692940682e+17, 1.27767692950682e+17, 1.27767692960682e+17, 1.27767692970682e+17, 1.27767692980682e+17, 1.27767692990682e+17, 1.27767693000682e+17, 1.277676930106821e+17, 1.27767693020682e+17, 1.27767693030682e+17, 1.27767693040682e+17, 1.27767693050682e+17, 1.27767693060682e+17, 1.27767693070682e+17, 1.27767693080682e+17, 1.27767693090682e+17, 1.27767693100682e+17, 1.27767693110682e+17, 1.27767693120682e+17, 1.27767693130682e+17, 1.27767693140682e+17, 1.27767693150682e+17, 1.27767693160682e+17, 1.27767693170682e+17, 1.27767693180682e+17, 1.27767693190682e+17, 1.27767693200682e+17, 1.27767693210682e+17, 1.27767693220682e+17, 1.27767693230682e+17, 1.27767693240682e+17, 1.27767693250682e+17, 1.27767693260682e+17, 1.277676932706821e+17, 1.27767693280682e+17, 1.27767693290682e+17, 1.27767693300682e+17, 1.27767693310682e+17, 1.27767693320682e+17, 1.27767693330682e+17, 1.27767693340682e+17, 1.27767693350682e+17, 1.27767693360682e+17, 1.27767693370682e+17, 1.27767693380682e+17, 1.27767693390682e+17, 1.27767693400682e+17, 1.27767693410682e+17, 1.27767693420682e+17, 1.27767693430682e+17, 1.27767693440682e+17, 1.27767693450682e+17, 1.27767693460682e+17, 1.27767693470682e+17, 1.27767693480682e+17, 1.27767693490682e+17, 1.27767693500682e+17, 1.27767693510682e+17, 1.27767693520682e+17, 1.277676935306821e+17, 1.27767693540682e+17, 1.27767693550682e+17, 1.27767693560682e+17, 1.27767693570682e+17, 1.27767693580682e+17, 1.27767693590682e+17, 1.27767693600682e+17, 1.27767693610682e+17, 1.27767693620682e+17, 1.27767693630682e+17, 1.27767693640682e+17, 1.27767693650682e+17, 1.27767693660682e+17, 1.27767693670682e+17, 1.27767693680682e+17, 1.27767693690682e+17, 1.27767693700682e+17, 1.27767693710682e+17, 1.27767693720682e+17, 1.27767693730682e+17, 1.27767693740682e+17, 1.27767693750682e+17, 1.27767693760682e+17, 1.27767693770682e+17, 1.27767693780682e+17, 1.27767693790682e+17, 1.27767693800682e+17, 1.27767693810682e+17, 1.27767693820682e+17, 1.27767693830682e+17, 1.27767693840682e+17, 1.27767693850682e+17, 1.27767693860682e+17, 1.27767693870682e+17, 1.27767693880682e+17, 1.27767693890682e+17, 1.27767693900682e+17, 1.27767693910682e+17, 1.27767693920682e+17, 1.27767693930682e+17, 1.27767693940682e+17, 1.27767693950682e+17, 1.27767693960682e+17, 1.27767693970682e+17, 1.27767693980682e+17, 1.27767693990682e+17, 1.27767694000682e+17, 1.27767694010682e+17, 1.27767694020682e+17, 1.27767694030682e+17, 1.27767694040682e+17, 1.27767694050682e+17, 1.27767694060682e+17, 1.27767694070682e+17, 1.27767694080682e+17, 1.27767694090682e+17, 1.27767694100682e+17, 1.27767694110682e+17, 1.27767694120682e+17, 1.27767694130682e+17, 1.27767694140682e+17, 1.27767694150682e+17, 1.277676941606821e+17, 1.27767694170682e+17, 1.27767694180682e+17, 1.27767694190682e+17, 1.27767694200682e+17, 1.27767694210682e+17, 1.27767694220682e+17, 1.27767694230682e+17, 1.27767694240682e+17, 1.27767694250682e+17, 1.27767694260682e+17, 1.27767694270682e+17, 1.27767694280682e+17, 1.27767694290682e+17, 1.27767694300682e+17, 1.27767694310682e+17, 1.27767694320682e+17, 1.27767694330682e+17, 1.27767694340682e+17, 1.27767694350682e+17, 1.27767694360682e+17, 1.27767694370682e+17, 1.27767694380682e+17, 1.27767694390682e+17, 1.27767694400682e+17, 1.27767694410682e+17, 1.277676944206821e+17, 1.27767694430682e+17, 1.27767694440682e+17, 1.27767694450682e+17, 1.27767694460682e+17, 1.27767694470682e+17, 1.27767694480682e+17},
			             {1.27767687110682e+17, 1.27767687120682e+17, 1.27767687130682e+17, 1.27767687140682e+17, 1.27767687150682e+17, 1.27767687160682e+17, 1.27767687170682e+17, 1.27767687180682e+17, 1.27767687190682e+17, 1.27767687200682e+17, 1.27767687210682e+17, 1.27767687220682e+17, 1.27767687230682e+17, 1.27767687240682e+17, 1.27767687250682e+17, 1.27767687260682e+17, 1.27767687270682e+17, 1.27767687280682e+17, 1.27767687290682e+17, 1.27767687300682e+17, 1.27767687310682e+17, 1.27767687320682e+17, 1.27767687330682e+17, 1.27767687340682e+17, 1.27767687350682e+17, 1.27767687360682e+17, 1.27767687370682e+17, 1.27767687380682e+17, 1.27767687390682e+17, 1.27767687400682e+17, 1.277676874106821e+17, 1.27767687420682e+17, 1.27767687430682e+17, 1.27767687440682e+17, 1.27767687450682e+17, 1.27767687460682e+17, 1.27767687470682e+17, 1.27767687480682e+17, 1.27767687490682e+17, 1.27767687500682e+17, 1.27767687510682e+17, 1.27767687520682e+17, 1.27767687530682e+17, 1.27767687540682e+17, 1.27767687550682e+17, 1.27767687560682e+17, 1.27767687570682e+17, 1.27767687580682e+17, 1.27767687590682e+17, 1.27767687600682e+17, 1.27767687610682e+17, 1.27767687620682e+17, 1.27767687630682e+17, 1.27767687640682e+17, 1.27767687650682e+17, 1.27767687660682e+17, 1.277676876706821e+17, 1.27767687680682e+17, 1.27767687690682e+17, 1.27767687700682e+17, 1.27767687710682e+17, 1.27767687720682e+17, 1.27767687730682e+17, 1.27767687740682e+17, 1.27767687750682e+17, 1.27767687760682e+17, 1.27767687770682e+17, 1.27767687780682e+17, 1.27767687790682e+17, 1.27767687800682e+17, 1.27767687810682e+17, 1.27767687820682e+17, 1.27767687830682e+17, 1.27767687840682e+17, 1.27767687850682e+17, 1.27767687860682e+17, 1.27767687870682e+17, 1.27767687880682e+17, 1.27767687890682e+17, 1.27767687900682e+17, 1.27767687910682e+17, 1.27767687920682e+17, 1.277676879306821e+17, 1.27767687940682e+17, 1.27767687950682e+17, 1.27767687960682e+17, 1.27767687970682e+17, 1.27767687980682e+17, 1.27767687990682e+17, 1.27767688000682e+17, 1.27767688010682e+17, 1.27767688020682e+17, 1.27767688030682e+17, 1.27767688040682e+17, 1.27767688050682e+17, 1.27767688060682e+17, 1.27767688070682e+17, 1.27767688080682e+17, 1.27767688090682e+17, 1.27767688100682e+17, 1.27767688110682e+17, 1.27767688120682e+17, 1.27767688130682e+17, 1.27767688140682e+17, 1.27767688150682e+17, 1.27767688160682e+17, 1.27767688170682e+17, 1.27767688180682e+17, 1.27767688190682e+17, 1.27767688200682e+17, 1.27767688210682e+17, 1.27767688220682e+17, 1.27767688230682e+17, 1.27767688240682e+17, 1.27767688250682e+17, 1.27767688260682e+17, 1.27767688270682e+17, 1.27767688280682e+17, 1.27767688290682e+17, 1.277676883006821e+17, 1.27767688310682e+17, 1.27767688320682e+17, 1.27767688330682e+17, 1.27767688340682e+17, 1.27767688350682e+17, 1.27767688360682e+17, 1.27767688370682e+17, 1.27767688380682e+17, 1.27767688390682e+17, 1.27767688400682e+17, 1.27767688410682e+17, 1.27767688420682e+17, 1.27767688430682e+17, 1.27767688440682e+17, 1.27767688450682e+17, 1.27767688460682e+17, 1.27767688470682e+17, 1.27767688480682e+17, 1.27767688490682e+17, 1.27767688500682e+17, 1.27767688510682e+17, 1.27767688520682e+17, 1.27767688530682e+17, 1.27767688540682e+17, 1.27767688550682e+17, 1.277676885606821e+17, 1.27767688570682e+17, 1.27767688580682e+17, 1.27767688590682e+17, 1.27767688600682e+17, 1.27767688610682e+17, 1.27767688620682e+17, 1.27767688630682e+17, 1.27767688640682e+17, 1.27767688650682e+17, 1.27767688660682e+17, 1.27767688670682e+17, 1.27767688680682e+17, 1.27767688690682e+17, 1.27767688700682e+17, 1.27767688710682e+17, 1.27767688720682e+17, 1.27767688730682e+17, 1.27767688740682e+17, 1.27767688750682e+17, 1.27767688760682e+17, 1.27767688770682e+17, 1.27767688780682e+17, 1.27767688790682e+17, 1.27767688800682e+17, 1.27767688810682e+17, 1.277676888206821e+17, 1.27767688830682e+17, 1.27767688840682e+17, 1.27767688850682e+17, 1.27767688860682e+17, 1.27767688870682e+17, 1.27767688880682e+17, 1.27767688890682e+17, 1.27767688900682e+17, 1.27767688910682e+17, 1.27767688920682e+17, 1.27767688930682e+17, 1.27767688940682e+17, 1.27767688950682e+17, 1.27767688960682e+17, 1.27767688970682e+17, 1.27767688980682e+17, 1.27767688990682e+17, 1.27767689000682e+17, 1.27767689010682e+17, 1.27767689020682e+17, 1.27767689030682e+17, 1.27767689040682e+17, 1.27767689050682e+17, 1.27767689060682e+17, 1.27767689070682e+17, 1.27767689080682e+17, 1.27767689090682e+17, 1.27767689100682e+17, 1.27767689110682e+17, 1.27767689120682e+17, 1.27767689130682e+17, 1.27767689140682e+17, 1.27767689150682e+17, 1.27767689160682e+17, 1.27767689170682e+17, 1.27767689180682e+17, 1.277676891906821e+17, 1.27767689200682e+17, 1.27767689210682e+17, 1.27767689220682e+17, 1.27767689230682e+17, 1.27767689240682e+17, 1.27767689250682e+17, 1.27767689260682e+17, 1.27767689270682e+17, 1.27767689280682e+17, 1.27767689290682e+17, 1.27767689300682e+17, 1.27767689310682e+17, 1.27767689320682e+17, 1.27767689330682e+17, 1.27767689340682e+17, 1.27767689350682e+17, 1.27767689360682e+17, 1.27767689370682e+17, 1.27767689380682e+17, 1.27767689390682e+17, 1.27767689400682e+17, 1.27767689410682e+17, 1.27767689420682e+17, 1.27767689430682e+17, 1.27767689440682e+17, 1.277676894506821e+17, 1.27767689460682e+17, 1.27767689470682e+17, 1.27767689480682e+17, 1.27767689490682e+17, 1.27767689500682e+17, 1.27767689510682e+17, 1.27767689520682e+17, 1.27767689530682e+17, 1.27767689540682e+17, 1.27767689550682e+17, 1.27767689560682e+17, 1.27767689570682e+17, 1.27767689580682e+17, 1.27767689590682e+17, 1.27767689600682e+17, 1.27767689610682e+17, 1.27767689620682e+17, 1.27767689630682e+17, 1.27767689640682e+17, 1.27767689650682e+17, 1.27767689660682e+17, 1.27767689670682e+17, 1.27767689680682e+17, 1.27767689690682e+17, 1.27767689700682e+17, 1.277676897106821e+17, 1.27767689720682e+17, 1.27767689730682e+17, 1.27767689740682e+17, 1.27767689750682e+17, 1.27767689760682e+17, 1.27767689770682e+17, 1.27767689780682e+17, 1.27767689790682e+17, 1.27767689800682e+17, 1.27767689810682e+17, 1.27767689820682e+17, 1.27767689830682e+17, 1.27767689840682e+17, 1.27767689850682e+17, 1.27767689860682e+17, 1.27767689870682e+17, 1.27767689880682e+17, 1.27767689890682e+17, 1.27767689900682e+17, 1.27767689910682e+17, 1.27767689920682e+17, 1.27767689930682e+17, 1.27767689940682e+17, 1.27767689950682e+17, 1.27767689960682e+17, 1.27767689970682e+17, 1.27767689980682e+17, 1.27767689990682e+17, 1.27767690000682e+17, 1.27767690010682e+17, 1.27767690020682e+17, 1.27767690030682e+17, 1.27767690040682e+17, 1.27767690050682e+17, 1.27767690060682e+17, 1.27767690070682e+17, 1.277676900806821e+17, 1.27767690090682e+17, 1.27767690100682e+17, 1.27767690110682e+17, 1.27767690120682e+17, 1.27767690130682e+17, 1.27767690140682e+17, 1.27767690150682e+17, 1.27767690160682e+17, 1.27767690170682e+17, 1.27767690180682e+17, 1.27767690190682e+17, 1.27767690200682e+17, 1.27767690210682e+17, 1.27767690220682e+17, 1.27767690230682e+17, 1.27767690240682e+17, 1.27767690250682e+17, 1.27767690260682e+17, 1.27767690270682e+17, 1.27767690280682e+17, 1.27767690290682e+17, 1.27767690300682e+17, 1.27767690310682e+17, 1.27767690320682e+17, 1.27767690330682e+17, 1.277676903406821e+17, 1.27767690350682e+17, 1.27767690360682e+17, 1.27767690370682e+17, 1.27767690380682e+17, 1.27767690390682e+17, 1.27767690400682e+17, 1.27767690410682e+17, 1.27767690420682e+17, 1.27767690430682e+17, 1.27767690440682e+17, 1.27767690450682e+17, 1.27767690460682e+17, 1.27767690470682e+17, 1.27767690480682e+17, 1.27767690490682e+17, 1.27767690500682e+17, 1.27767690510682e+17, 1.27767690520682e+17, 1.27767690530682e+17, 1.27767690540682e+17, 1.27767690550682e+17, 1.27767690560682e+17, 1.27767690570682e+17, 1.27767690580682e+17, 1.27767690590682e+17, 1.277676906006821e+17, 1.27767690610682e+17, 1.27767690620682e+17, 1.27767690630682e+17, 1.27767690640682e+17, 1.27767690650682e+17, 1.27767690660682e+17, 1.27767690670682e+17, 1.27767690680682e+17, 1.27767690690682e+17, 1.27767690700682e+17, 1.27767690710682e+17, 1.27767690720682e+17, 1.27767690730682e+17, 1.27767690740682e+17, 1.27767690750682e+17, 1.27767690760682e+17, 1.27767690770682e+17, 1.27767690780682e+17, 1.27767690790682e+17, 1.27767690800682e+17, 1.27767690810682e+17, 1.27767690820682e+17, 1.27767690830682e+17, 1.27767690840682e+17, 1.27767690850682e+17, 1.27767690860682e+17, 1.27767690870682e+17, 1.27767690880682e+17, 1.27767690890682e+17, 1.27767690900682e+17, 1.27767690910682e+17, 1.27767690920682e+17, 1.27767690930682e+17, 1.27767690940682e+17, 1.27767690950682e+17, 1.27767690960682e+17, 1.27767690970682e+17, 1.27767690980682e+17, 1.27767690990682e+17, 1.27767691000682e+17, 1.27767691010682e+17, 1.27767691020682e+17, 1.27767691030682e+17, 1.27767691040682e+17, 1.27767691050682e+17, 1.27767691060682e+17, 1.27767691070682e+17, 1.27767691080682e+17, 1.27767691090682e+17, 1.27767691100682e+17, 1.27767691110682e+17, 1.27767691120682e+17, 1.27767691130682e+17, 1.27767691140682e+17, 1.27767691150682e+17, 1.27767691160682e+17, 1.27767691170682e+17, 1.27767691180682e+17, 1.27767691190682e+17, 1.27767691200682e+17, 1.27767691210682e+17, 1.27767691220682e+17, 1.277676912306821e+17, 1.27767691240682e+17, 1.27767691250682e+17, 1.27767691260682e+17, 1.27767691270682e+17, 1.27767691280682e+17, 1.27767691290682e+17, 1.27767691300682e+17, 1.27767691310682e+17, 1.27767691320682e+17, 1.27767691330682e+17, 1.27767691340682e+17, 1.27767691350682e+17, 1.27767691360682e+17, 1.27767691370682e+17, 1.27767691380682e+17, 1.27767691390682e+17, 1.27767691400682e+17, 1.27767691410682e+17, 1.27767691420682e+17, 1.27767691430682e+17, 1.27767691440682e+17, 1.27767691450682e+17, 1.27767691460682e+17},
			             {1.27767706080682e+17, 1.27767706090682e+17, 1.27767706100682e+17, 1.27767706110682e+17, 1.27767706120682e+17, 1.27767706130682e+17, 1.277677061406821e+17, 1.27767706150682e+17, 1.27767706160682e+17, 1.27767706170682e+17, 1.27767706180682e+17, 1.27767706190682e+17, 1.27767706200682e+17, 1.27767706210682e+17},
			             {1.27767702330682e+17, 1.27767702340682e+17, 1.27767702350682e+17, 1.27767702360682e+17, 1.27767702370682e+17, 1.27767702380682e+17, 1.27767702390682e+17, 1.27767702400682e+17, 1.27767702410682e+17, 1.27767702420682e+17, 1.27767702430682e+17},
			             {1.27767702600682e+17, 1.27767702610682e+17, 1.27767702620682e+17, 1.27767702630682e+17, 1.27767702640682e+17},
			             {1.27767703200682e+17, 1.277677032106821e+17, 1.27767703220682e+17, 1.27767703230682e+17, 1.27767703240682e+17},
			             {1.27767703100682e+17, 1.27767703110682e+17, 1.27767703120682e+17, 1.27767703130682e+17, 1.27767703140682e+17, 1.27767703150682e+17, 1.27767703160682e+17},
			             {1.27767707040682e+17, 1.27767707050682e+17, 1.27767707060682e+17, 1.27767707070682e+17, 1.27767707080682e+17, 1.27767707090682e+17, 1.27767707100682e+17, 1.27767707110682e+17, 1.27767707120682e+17, 1.27767707130682e+17, 1.27767707140682e+17, 1.27767707150682e+17, 1.27767707160682e+17, 1.27767707170682e+17, 1.27767707180682e+17, 1.27767707190682e+17, 1.27767707200682e+17, 1.27767707210682e+17, 1.27767707220682e+17, 1.27767707230682e+17, 1.27767707240682e+17, 1.27767707250682e+17, 1.27767707260682e+17, 1.27767707270682e+17, 1.27767707280682e+17, 1.27767707290682e+17, 1.27767707300682e+17, 1.27767707310682e+17, 1.27767707320682e+17, 1.27767707330682e+17, 1.27767707340682e+17, 1.27767707350682e+17, 1.27767707360682e+17, 1.27767707370682e+17, 1.27767707380682e+17, 1.27767707390682e+17, 1.27767707400682e+17, 1.27767707410682e+17, 1.27767707420682e+17, 1.27767707430682e+17, 1.27767707440682e+17, 1.27767707450682e+17, 1.27767707460682e+17, 1.27767707470682e+17, 1.27767707480682e+17, 1.27767707490682e+17, 1.27767707500682e+17, 1.27767707510682e+17, 1.27767707520682e+17, 1.27767707530682e+17, 1.27767707540682e+17, 1.27767707550682e+17, 1.27767707560682e+17, 1.27767707570682e+17, 1.27767707580682e+17, 1.27767707590682e+17, 1.27767707600682e+17, 1.27767707610682e+17, 1.27767707620682e+17, 1.27767707630682e+17, 1.27767707640682e+17, 1.27767707650682e+17, 1.277677076606821e+17, 1.27767707670682e+17, 1.27767707680682e+17, 1.27767707690682e+17, 1.27767707700682e+17, 1.27767707710682e+17, 1.27767707720682e+17, 1.27767707730682e+17, 1.27767707740682e+17, 1.27767707750682e+17, 1.27767707760682e+17, 1.27767707770682e+17, 1.27767707780682e+17, 1.27767707790682e+17, 1.27767707800682e+17, 1.27767707810682e+17, 1.27767707820682e+17, 1.27767707830682e+17, 1.27767707840682e+17, 1.27767707850682e+17, 1.27767707860682e+17, 1.27767707870682e+17, 1.27767707880682e+17, 1.27767707890682e+17, 1.27767707900682e+17, 1.27767707910682e+17, 1.277677079206821e+17, 1.27767707930682e+17, 1.27767707940682e+17, 1.27767707950682e+17, 1.27767707960682e+17, 1.27767707970682e+17, 1.27767707980682e+17, 1.27767707990682e+17, 1.27767708000682e+17, 1.27767708010682e+17, 1.27767708020682e+17, 1.27767708030682e+17, 1.27767708040682e+17, 1.27767708050682e+17, 1.27767708060682e+17, 1.27767708070682e+17, 1.27767708080682e+17, 1.27767708090682e+17, 1.27767708100682e+17, 1.27767708110682e+17, 1.27767708120682e+17, 1.27767708130682e+17, 1.27767708140682e+17, 1.27767708150682e+17, 1.27767708160682e+17, 1.27767708170682e+17, 1.277677081806821e+17, 1.27767708190682e+17, 1.27767708200682e+17, 1.27767708210682e+17, 1.27767708220682e+17, 1.27767708230682e+17, 1.27767708240682e+17, 1.27767708250682e+17, 1.27767708260682e+17, 1.27767708270682e+17, 1.27767708280682e+17, 1.27767708290682e+17, 1.27767708300682e+17, 1.27767708310682e+17, 1.27767708320682e+17, 1.27767708330682e+17, 1.27767708340682e+17, 1.27767708350682e+17, 1.27767708360682e+17, 1.27767708370682e+17, 1.27767708380682e+17, 1.27767708390682e+17, 1.27767708400682e+17, 1.27767708410682e+17, 1.27767708420682e+17, 1.27767708430682e+17, 1.27767708440682e+17, 1.27767708450682e+17, 1.27767708460682e+17, 1.27767708470682e+17, 1.27767708480682e+17, 1.27767708490682e+17, 1.27767708500682e+17, 1.27767708510682e+17, 1.27767708520682e+17, 1.27767708530682e+17, 1.27767708540682e+17, 1.277677085506821e+17, 1.27767708560682e+17, 1.27767708570682e+17, 1.27767708580682e+17, 1.27767708590682e+17, 1.27767708600682e+17, 1.27767708610682e+17, 1.27767708620682e+17, 1.27767708630682e+17, 1.27767708640682e+17, 1.27767708650682e+17, 1.27767708660682e+17, 1.27767708670682e+17, 1.27767708680682e+17, 1.27767708690682e+17, 1.27767708700682e+17, 1.27767708710682e+17, 1.27767708720682e+17, 1.27767708730682e+17, 1.27767708740682e+17, 1.27767708750682e+17, 1.27767708760682e+17, 1.27767708770682e+17, 1.27767708780682e+17, 1.27767708790682e+17, 1.27767708800682e+17, 1.277677088106821e+17, 1.27767708820682e+17, 1.27767708830682e+17, 1.27767708840682e+17, 1.27767708850682e+17, 1.27767708860682e+17, 1.27767708870682e+17, 1.27767708880682e+17, 1.27767708890682e+17, 1.27767708900682e+17, 1.27767708910682e+17, 1.27767708920682e+17, 1.27767708930682e+17, 1.27767708940682e+17, 1.27767708950682e+17, 1.27767708960682e+17, 1.27767708970682e+17, 1.27767708980682e+17, 1.27767708990682e+17, 1.27767709000682e+17, 1.27767709010682e+17, 1.27767709020682e+17, 1.27767709030682e+17, 1.27767709040682e+17, 1.27767709050682e+17, 1.27767709060682e+17, 1.277677090706821e+17, 1.27767709080682e+17, 1.27767709090682e+17, 1.27767709100682e+17, 1.27767709110682e+17, 1.27767709120682e+17, 1.27767709130682e+17, 1.27767709140682e+17, 1.27767709150682e+17, 1.27767709160682e+17, 1.27767709170682e+17, 1.27767709180682e+17, 1.27767709190682e+17, 1.27767709200682e+17, 1.27767709210682e+17, 1.27767709220682e+17, 1.27767709230682e+17, 1.27767709240682e+17, 1.27767709250682e+17, 1.27767709260682e+17, 1.27767709270682e+17, 1.27767709280682e+17, 1.27767709290682e+17, 1.27767709300682e+17, 1.27767709310682e+17, 1.27767709320682e+17, 1.27767709330682e+17, 1.27767709340682e+17, 1.27767709350682e+17, 1.27767709360682e+17, 1.27767709370682e+17, 1.27767709380682e+17, 1.27767709390682e+17, 1.27767709420682e+17, 1.27767709430682e+17, 1.277677094406821e+17, 1.27767709450682e+17, 1.27767709460682e+17, 1.27767709470682e+17, 1.27767709480682e+17, 1.27767709490682e+17, 1.27767709500682e+17, 1.27767709510682e+17, 1.27767709520682e+17, 1.27767709530682e+17, 1.27767709540682e+17, 1.27767709550682e+17, 1.27767709560682e+17, 1.27767709570682e+17, 1.27767709580682e+17, 1.27767709590682e+17, 1.27767709600682e+17, 1.27767709610682e+17, 1.27767709620682e+17, 1.27767709630682e+17, 1.27767709640682e+17, 1.27767709650682e+17, 1.27767709660682e+17, 1.27767709670682e+17, 1.27767709680682e+17, 1.27767709690682e+17, 1.277677097006821e+17, 1.27767709710682e+17, 1.27767709720682e+17, 1.27767709730682e+17, 1.27767709740682e+17, 1.27767709750682e+17, 1.27767709760682e+17, 1.27767709770682e+17, 1.27767709780682e+17, 1.27767709790682e+17, 1.27767709800682e+17, 1.27767709810682e+17, 1.27767709820682e+17, 1.27767709830682e+17, 1.27767709840682e+17, 1.27767709850682e+17, 1.27767709860682e+17, 1.27767709870682e+17, 1.27767709880682e+17, 1.27767709890682e+17, 1.27767709900682e+17, 1.27767709910682e+17, 1.27767709920682e+17, 1.27767709930682e+17, 1.27767709940682e+17, 1.27767709950682e+17, 1.277677099606821e+17, 1.27767709970682e+17, 1.27767709980682e+17, 1.27767709990682e+17, 1.27767710000682e+17, 1.27767710010682e+17, 1.27767710020682e+17, 1.27767710030682e+17, 1.27767710040682e+17, 1.27767710050682e+17, 1.27767710060682e+17, 1.27767710070682e+17, 1.27767710080682e+17, 1.27767710090682e+17, 1.27767710100682e+17, 1.27767710110682e+17, 1.27767710120682e+17, 1.27767710130682e+17, 1.27767710140682e+17, 1.27767710150682e+17, 1.27767710160682e+17, 1.27767710170682e+17, 1.27767710180682e+17, 1.27767710190682e+17, 1.27767710200682e+17, 1.27767710210682e+17, 1.27767710220682e+17, 1.27767710230682e+17, 1.27767710240682e+17, 1.27767710250682e+17, 1.27767710260682e+17, 1.27767710270682e+17, 1.27767710280682e+17, 1.27767710290682e+17, 1.27767710300682e+17, 1.27767710310682e+17, 1.27767710320682e+17, 1.277677103306821e+17, 1.27767710340682e+17, 1.27767710350682e+17, 1.27767710360682e+17, 1.27767710370682e+17, 1.27767710380682e+17, 1.27767710390682e+17, 1.27767710400682e+17, 1.27767710410682e+17, 1.27767710420682e+17, 1.27767710430682e+17, 1.27767710440682e+17, 1.27767710450682e+17, 1.27767710460682e+17, 1.27767710470682e+17, 1.27767710480682e+17, 1.27767710490682e+17, 1.27767710500682e+17, 1.27767710510682e+17, 1.27767710520682e+17, 1.27767710530682e+17, 1.27767710540682e+17, 1.27767710550682e+17, 1.27767710560682e+17, 1.27767710570682e+17, 1.27767710580682e+17, 1.277677105906821e+17, 1.27767710600682e+17, 1.27767710610682e+17, 1.27767710620682e+17, 1.27767710630682e+17, 1.27767710640682e+17, 1.27767710650682e+17, 1.27767710660682e+17, 1.27767710670682e+17, 1.27767710680682e+17, 1.27767710690682e+17, 1.27767710700682e+17, 1.27767710710682e+17, 1.27767710720682e+17, 1.27767710730682e+17, 1.27767710740682e+17, 1.27767710750682e+17, 1.27767710760682e+17, 1.27767710770682e+17, 1.27767710780682e+17, 1.27767710790682e+17, 1.27767710800682e+17, 1.27767710810682e+17, 1.27767710820682e+17, 1.27767710830682e+17, 1.27767710840682e+17, 1.277677108506821e+17, 1.27767710860682e+17, 1.277677108678696e+17, 1.27767710880682e+17, 1.277677108903695e+17, 1.277677108975571e+17, 1.27767710910682e+17, 1.27767710920682e+17, 1.277677109297445e+17, 1.277677109359945e+17, 1.27767710950682e+17, 1.27767710960682e+17, 1.27767710970682e+17, 1.27767710980682e+17, 1.27767710990682e+17, 1.27767711000682e+17, 1.277677110070883e+17, 1.277677110167757e+17, 1.27767711030682e+17, 1.27767711040682e+17, 1.27767711050682e+17, 1.27767711060682e+17, 1.277677110699008e+17, 1.27767711080682e+17, 1.27767711090682e+17, 1.27767711100682e+17, 1.27767711110682e+17, 1.277677111202132e+17, 1.27767711130682e+17, 1.27767711140682e+17, 1.27767711150682e+17, 1.27767711160682e+17, 1.27767711170057e+17, 1.27767711180682e+17, 1.27767711190682e+17, 1.27767711200682e+17, 1.27767711210682e+17, 1.277677112202132e+17, 1.27767711230682e+17, 1.27767711240682e+17, 1.27767711250682e+17, 1.27767711260682e+17, 1.277677112694319e+17, 1.27767711280682e+17, 1.27767711290682e+17, 1.27767711300682e+17, 1.27767711310682e+17, 1.277677113195882e+17, 1.27767711330682e+17, 1.27767711340682e+17, 1.27767711350682e+17, 1.27767711360682e+17, 1.27767711370682e+17, 1.277677113803695e+17, 1.27767711390682e+17, 1.27767711400682e+17, 1.27767711410682e+17, 1.27767711420682e+17, 1.277677114295882e+17, 1.27767711440682e+17, 1.27767711450682e+17, 1.27767711460682e+17, 1.27767711470682e+17, 1.277677114792756e+17, 1.27767711490682e+17, 1.27767711500682e+17, 1.27767711510682e+17, 1.27767711520682e+17, 1.277677115295882e+17, 1.27767711540682e+17, 1.27767711550682e+17, 1.27767711560682e+17, 1.27767711570682e+17, 1.277677115797445e+17, 1.27767711590682e+17, 1.27767711600682e+17, 1.27767711610682e+17, 1.27767711620682e+17, 1.277677116295884e+17, 1.27767711640682e+17, 1.27767711650682e+17, 1.27767711660682e+17, 1.27767711670682e+17, 1.277677116799008e+17, 1.27767711690682e+17, 1.27767711700682e+17, 1.27767711710682e+17, 1.27767711720682e+17, 1.27767711730057e+17, 1.277677117406821e+17, 1.27767711750682e+17, 1.27767711760682e+17, 1.27767711770682e+17, 1.277677117799007e+17, 1.27767711790682e+17, 1.27767711800682e+17, 1.27767711810682e+17, 1.27767711820682e+17, 1.277677118302132e+17, 1.27767711840682e+17, 1.27767711850682e+17, 1.27767711860682e+17, 1.27767711870682e+17, 1.277677118792758e+17, 1.27767711890682e+17, 1.27767711900682e+17, 1.27767711910682e+17, 1.27767711920682e+17, 1.27767711930682e+17, 1.27767711940682e+17, 1.27767711950682e+17, 1.27767711960682e+17, 1.27767711970682e+17, 1.277677119803695e+17, 1.277677119903695e+17, 1.277677120006821e+17, 1.27767712010682e+17, 1.27767712020682e+17, 1.27767712030682e+17, 1.277677120395884e+17, 1.27767712050682e+17, 1.27767712060682e+17, 1.27767712070682e+17, 1.27767712080682e+17, 1.277677120902132e+17, 1.27767712100682e+17, 1.27767712110682e+17, 1.27767712120682e+17, 1.27767712130682e+17, 1.277677121402132e+17, 1.27767712150682e+17, 1.27767712160682e+17, 1.27767712170682e+17, 1.27767712180682e+17, 1.277677121895882e+17, 1.27767712200682e+17, 1.27767712210682e+17, 1.27767712220682e+17, 1.27767712230682e+17, 1.277677122397445e+17, 1.27767712250682e+17, 1.27767712260682e+17, 1.27767712270682e+17, 1.27767712280682e+17, 1.277677122899008e+17, 1.27767712300682e+17, 1.27767712310682e+17, 1.27767712320682e+17, 1.27767712330682e+17, 1.277677123397445e+17, 1.27767712350682e+17, 1.27767712360682e+17, 1.277677123706821e+17, 1.27767712380682e+17, 1.27767712390057e+17, 1.27767712400682e+17, 1.27767712410682e+17, 1.27767712420682e+17, 1.27767712430682e+17, 1.277677124397444e+17, 1.27767712450682e+17, 1.27767712460682e+17, 1.27767712470682e+17, 1.277677124799007e+17, 1.27767712490682e+17, 1.27767712500682e+17, 1.27767712510682e+17, 1.27767712520057e+17, 1.27767712530682e+17, 1.27767712540682e+17, 1.27767712550682e+17, 1.27767712560057e+17, 1.27767712570682e+17, 1.27767712580682e+17, 1.27767712590682e+17, 1.277677126002132e+17, 1.27767712610682e+17, 1.27767712620682e+17, 1.277677126306821e+17, 1.277677126394319e+17, 1.27767712650682e+17, 1.27767712660682e+17, 1.27767712670682e+17, 1.277677126794319e+17, 1.27767712690682e+17, 1.27767712700682e+17, 1.27767712710682e+17, 1.277677127202132e+17, 1.27767712730682e+17, 1.27767712740682e+17, 1.27767712750682e+17, 1.277677127594321e+17, 1.27767712770682e+17, 1.27767712780682e+17, 1.27767712790682e+17, 1.277677127995884e+17, 1.27767712810682e+17, 1.27767712820682e+17, 1.27767712830682e+17, 1.277677128397445e+17, 1.27767712850682e+17, 1.27767712860682e+17, 1.27767712870682e+17, 1.277677128795882e+17, 1.277677128906821e+17, 1.27767712900682e+17, 1.27767712910682e+17, 1.277677129195882e+17, 1.27767712930682e+17, 1.27767712940682e+17, 1.27767712950682e+17, 1.277677129597444e+17, 1.27767712970682e+17, 1.27767712980682e+17, 1.27767712990682e+17, 1.277677129999007e+17, 1.27767713010682e+17, 1.27767713020682e+17, 1.27767713030682e+17, 1.277677130397445e+17, 1.27767713050682e+17, 1.27767713060682e+17, 1.27767713070682e+17, 1.277677130799008e+17, 1.27767713090682e+17, 1.27767713100682e+17, 1.27767713110682e+17, 1.277677131199008e+17, 1.27767713130682e+17, 1.27767713140682e+17, 1.27767713150682e+17, 1.27767713160057e+17, 1.27767713170682e+17, 1.27767713180682e+17, 1.27767713190682e+17, 1.277677131992758e+17, 1.27767713210682e+17, 1.27767713220682e+17, 1.27767713230682e+17, 1.277677132400571e+17, 1.27767713250682e+17, 1.277677132606821e+17, 1.27767713270682e+17, 1.277677132802132e+17, 1.27767713290682e+17, 1.27767713300682e+17, 1.27767713310682e+17, 1.277677133192758e+17, 1.27767713330682e+17, 1.27767713340682e+17, 1.27767713350682e+17, 1.277677133595882e+17, 1.27767713370682e+17, 1.27767713380682e+17, 1.27767713390682e+17, 1.277677133994319e+17, 1.27767713410682e+17, 1.27767713420682e+17, 1.27767713430682e+17, 1.277677134394321e+17, 1.27767713450682e+17, 1.27767713460682e+17, 1.27767713470682e+17, 1.277677134795882e+17, 1.27767713490682e+17, 1.27767713500682e+17, 1.27767713510682e+17, 1.277677135202132e+17, 1.27767713530682e+17, 1.27767713540682e+17, 1.27767713550682e+17, 1.277677135595884e+17, 1.27767713570682e+17, 1.27767713580682e+17, 1.27767713590682e+17, 1.277677135995882e+17, 1.27767713610682e+17, 1.27767713620682e+17, 1.27767713630682e+17, 1.277677136397445e+17, 1.27767713650682e+17, 1.27767713660682e+17, 1.27767713670682e+17, 1.277677136799008e+17, 1.27767713690682e+17, 1.27767713700682e+17, 1.27767713710682e+17, 1.277677137197445e+17, 1.27767713730682e+17, 1.27767713740682e+17, 1.27767713750682e+17, 1.277677137599007e+17, 1.27767713770682e+17, 1.277677137806821e+17, 1.27767713790682e+17, 1.27767713800057e+17, 1.27767713810682e+17, 1.27767713820682e+17, 1.27767713830682e+17, 1.277677138402132e+17, 1.27767713850682e+17, 1.27767713860682e+17, 1.27767713870682e+17, 1.27767713880057e+17, 1.27767713890682e+17, 1.27767713900682e+17, 1.27767713910682e+17, 1.277677139202132e+17, 1.27767713930682e+17, 1.27767713940682e+17, 1.27767713950682e+17, 1.277677139592758e+17, 1.27767713970682e+17, 1.27767713980682e+17, 1.27767713990682e+17, 1.277677139994321e+17, 1.27767714010682e+17, 1.27767714020682e+17, 1.27767714030682e+17, 1.277677140402132e+17, 1.27767714050682e+17, 1.27767714060682e+17, 1.27767714070682e+17, 1.277677140794319e+17, 1.27767714090682e+17, 1.27767714100682e+17, 1.27767714110682e+17, 1.27767714120057e+17, 1.27767714130682e+17, 1.27767714140682e+17, 1.27767714150682e+17, 1.277677141602132e+17, 1.27767714170682e+17, 1.27767714180682e+17, 1.27767714190682e+17, 1.277677141994319e+17, 1.27767714210682e+17, 1.27767714220682e+17, 1.27767714230682e+17, 1.277677142395882e+17, 1.27767714250682e+17, 1.27767714260682e+17, 1.27767714270682e+17, 1.277677142797445e+17, 1.27767714290682e+17, 1.27767714300682e+17, 1.27767714310682e+17, 1.277677143199008e+17, 1.27767714330682e+17, 1.27767714340682e+17, 1.27767714350682e+17, 1.277677143594319e+17, 1.27767714370682e+17, 1.27767714380682e+17, 1.27767714390682e+17, 1.277677143997445e+17, 1.277677144106821e+17, 1.27767714420682e+17, 1.27767714430682e+17, 1.277677144399008e+17, 1.27767714450682e+17, 1.27767714460682e+17, 1.27767714470682e+17, 1.277677144800571e+17, 1.27767714490682e+17, 1.27767714500682e+17, 1.27767714510682e+17, 1.277677145194321e+17, 1.27767714530682e+17, 1.27767714540682e+17, 1.27767714550682e+17, 1.27767714560057e+17, 1.27767714570682e+17, 1.27767714580682e+17, 1.27767714590682e+17, 1.277677146002132e+17, 1.27767714610682e+17, 1.27767714620682e+17, 1.27767714630682e+17, 1.277677146392758e+17, 1.27767714650682e+17, 1.27767714660682e+17, 1.277677146706821e+17, 1.277677146794319e+17, 1.27767714690682e+17, 1.27767714700682e+17, 1.27767714710682e+17, 1.277677147202132e+17, 1.27767714730682e+17, 1.27767714740682e+17, 1.27767714750682e+17, 1.277677147592758e+17, 1.27767714770682e+17, 1.27767714780682e+17, 1.27767714790682e+17, 1.277677147994321e+17, 1.27767714810682e+17, 1.27767714820682e+17, 1.27767714830682e+17, 1.277677148395884e+17, 1.27767714850682e+17, 1.27767714860682e+17, 1.27767714870682e+17, 1.277677148794319e+17, 1.27767714890682e+17, 1.27767714900682e+17, 1.27767714910682e+17, 1.277677149195882e+17, 1.277677149306821e+17, 1.27767714940682e+17, 1.277677149486508e+17, 1.277677149586508e+17, 1.27767714970682e+17, 1.27767714980682e+17, 1.27767714990682e+17, 1.277677149999008e+17, 1.27767715010682e+17, 1.27767715020682e+17, 1.27767715030682e+17, 1.277677150395884e+17, 1.27767715050682e+17, 1.27767715060682e+17, 1.27767715070682e+17, 1.277677150797445e+17, 1.27767715090682e+17, 1.27767715100682e+17, 1.27767715110682e+17, 1.277677151199008e+17, 1.27767715130682e+17, 1.27767715140682e+17, 1.27767715150682e+17, 1.27767715160057e+17, 1.27767715170682e+17, 1.27767715180682e+17, 1.27767715190682e+17, 1.277677151999008e+17, 1.27767715210682e+17, 1.27767715220682e+17, 1.27767715230682e+17, 1.277677152399008e+17, 1.27767715250682e+17, 1.27767715260682e+17, 1.27767715270682e+17, 1.277677152799007e+17, 1.27767715290682e+17, 1.277677153006821e+17, 1.27767715310682e+17, 1.27767715320057e+17, 1.27767715330682e+17, 1.27767715340682e+17, 1.27767715350682e+17, 1.277677153602132e+17, 1.27767715370682e+17, 1.27767715380682e+17, 1.27767715390682e+17, 1.277677153992758e+17, 1.27767715410682e+17, 1.27767715420682e+17, 1.27767715430682e+17, 1.277677154394319e+17, 1.27767715450682e+17, 1.27767715460682e+17, 1.27767715470682e+17, 1.277677154800571e+17, 1.27767715490682e+17, 1.27767715500682e+17, 1.27767715510682e+17, 1.277677155194321e+17, 1.27767715530682e+17, 1.27767715540682e+17, 1.27767715550682e+17, 1.277677155595884e+17, 1.27767715570682e+17, 1.27767715580682e+17, 1.27767715590682e+17, 1.277677155997445e+17, 1.27767715610682e+17, 1.27767715620682e+17, 1.27767715630682e+17, 1.277677156397445e+17, 1.27767715650682e+17, 1.27767715660682e+17, 1.27767715670682e+17, 1.277677156795882e+17, 1.27767715690682e+17, 1.27767715700682e+17, 1.27767715710682e+17, 1.277677157197445e+17, 1.27767715730682e+17, 1.27767715740682e+17, 1.27767715750682e+17, 1.277677157599008e+17, 1.27767715770682e+17, 1.27767715780682e+17, 1.27767715790682e+17, 1.27767715800682e+17, 1.27767715810682e+17, 1.277677158206821e+17, 1.27767715830682e+17, 1.277677158399008e+17, 1.27767715850682e+17, 1.27767715860682e+17, 1.27767715870682e+17, 1.27767715880057e+17, 1.27767715890682e+17, 1.27767715900682e+17, 1.27767715910682e+17, 1.277677159202132e+17, 1.27767715930682e+17, 1.27767715940682e+17, 1.27767715950682e+17, 1.277677159597445e+17, 1.27767715970682e+17, 1.27767715980682e+17, 1.27767715990682e+17, 1.277677160000571e+17, 1.27767716010682e+17, 1.27767716020682e+17, 1.27767716030682e+17, 1.277677160402132e+17, 1.27767716050682e+17, 1.27767716060682e+17, 1.27767716070682e+17, 1.277677160794321e+17, 1.27767716090682e+17, 1.27767716100682e+17, 1.27767716110682e+17, 1.277677161195884e+17, 1.27767716130682e+17, 1.27767716140682e+17, 1.27767716150682e+17, 1.277677161592758e+17, 1.27767716170682e+17, 1.27767716180682e+17, 1.277677161906821e+17, 1.277677161994319e+17, 1.27767716210682e+17, 1.27767716220682e+17, 1.27767716230682e+17, 1.277677162395882e+17, 1.27767716250682e+17, 1.27767716260682e+17, 1.27767716270682e+17, 1.277677162797445e+17, 1.27767716290682e+17, 1.27767716300682e+17, 1.27767716310682e+17, 1.277677163203695e+17, 1.27767716330682e+17, 1.27767716340682e+17, 1.27767716350682e+17, 1.277677163595882e+17, 1.27767716370682e+17, 1.27767716380682e+17, 1.27767716390682e+17, 1.277677164005257e+17, 1.27767716410682e+17, 1.27767716420682e+17, 1.27767716430682e+17, 1.277677164399008e+17, 1.277677164506821e+17, 1.27767716460682e+17, 1.27767716470682e+17, 1.277677164799008e+17, 1.27767716490682e+17, 1.27767716500682e+17, 1.27767716510682e+17, 1.277677165200571e+17, 1.27767716530682e+17, 1.27767716540682e+17, 1.27767716550682e+17, 1.277677165597445e+17, 1.27767716570682e+17, 1.27767716580682e+17, 1.27767716590682e+17, 1.27767716600057e+17, 1.27767716610682e+17, 1.27767716620682e+17, 1.27767716630682e+17, 1.277677166402132e+17, 1.27767716650682e+17, 1.27767716660682e+17, 1.27767716670682e+17, 1.277677166792758e+17, 1.27767716690682e+17, 1.27767716700682e+17, 1.277677167106821e+17, 1.277677167194319e+17, 1.27767716730682e+17, 1.27767716740682e+17, 1.27767716750682e+17, 1.277677167602132e+17, 1.27767716770682e+17, 1.27767716780682e+17, 1.27767716790682e+17, 1.277677167992758e+17, 1.27767716810682e+17, 1.27767716820682e+17, 1.27767716830682e+17, 1.277677168394321e+17, 1.27767716850682e+17, 1.27767716860682e+17, 1.27767716870682e+17, 1.277677168795884e+17, 1.27767716890682e+17, 1.27767716900682e+17, 1.27767716910682e+17, 1.277677169202132e+17, 1.27767716930682e+17, 1.27767716940682e+17, 1.27767716950682e+17, 1.277677169594319e+17, 1.27767716970682e+17, 1.27767716980682e+17, 1.27767716990682e+17, 1.277677169995882e+17, 1.27767717010682e+17, 1.27767717020682e+17, 1.27767717030682e+17, 1.277677170397444e+17, 1.27767717050682e+17, 1.27767717060682e+17, 1.27767717070682e+17, 1.277677170794321e+17, 1.27767717090682e+17, 1.27767717100682e+17, 1.27767717110682e+17, 1.277677171197445e+17, 1.27767717130682e+17, 1.27767717140682e+17, 1.27767717150682e+17, 1.277677171599008e+17, 1.27767717170682e+17, 1.27767717180682e+17, 1.27767717190682e+17, 1.27767717200057e+17, 1.27767717210682e+17, 1.27767717220682e+17, 1.27767717230682e+17, 1.27767717240057e+17, 1.27767717250682e+17, 1.27767717260682e+17, 1.27767717270682e+17, 1.277677172797445e+17, 1.27767717290682e+17, 1.27767717300682e+17, 1.27767717310682e+17, 1.277677173200571e+17, 1.27767717330682e+17, 1.277677173406821e+17, 1.27767717350682e+17, 1.277677173602132e+17, 1.27767717370682e+17, 1.27767717380682e+17, 1.27767717390682e+17, 1.277677173992758e+17, 1.27767717410682e+17, 1.27767717420682e+17, 1.27767717430682e+17, 1.27767717440057e+17, 1.27767717450682e+17, 1.27767717460682e+17, 1.27767717470682e+17, 1.277677174802131e+17, 1.27767717490682e+17, 1.27767717500682e+17, 1.27767717510682e+17, 1.277677175194321e+17, 1.27767717530682e+17, 1.27767717540682e+17, 1.27767717550682e+17, 1.277677175602132e+17, 1.27767717570682e+17, 1.27767717580682e+17, 1.27767717590682e+17, 1.277677176002132e+17, 1.27767717610682e+17, 1.27767717620682e+17, 1.27767717630682e+17, 1.277677176392756e+17, 1.27767717650682e+17, 1.27767717660682e+17, 1.27767717670682e+17, 1.277677176795882e+17, 1.27767717690682e+17, 1.27767717700682e+17, 1.27767717710682e+17, 1.277677177197445e+17, 1.27767717730682e+17, 1.27767717740682e+17, 1.27767717750682e+17, 1.277677177599008e+17, 1.27767717770682e+17, 1.27767717780682e+17, 1.27767717790682e+17, 1.277677177999008e+17, 1.27767717810682e+17, 1.27767717820682e+17, 1.27767717830682e+17, 1.277677178397445e+17, 1.27767717850682e+17, 1.27767717860682e+17, 1.27767717870682e+17, 1.277677178799008e+17, 1.27767717890682e+17, 1.27767717900682e+17, 1.27767717910682e+17, 1.27767717920057e+17, 1.27767717930682e+17, 1.27767717940682e+17, 1.27767717950682e+17, 1.27767717960682e+17, 1.27767717970682e+17, 1.27767717980682e+17, 1.27767717990682e+17, 1.27767718000682e+17, 1.27767718010682e+17, 1.27767718020682e+17, 1.27767718030682e+17, 1.277677180391195e+17, 1.277677180480257e+17, 1.27767718060682e+17, 1.27767718070682e+17, 1.27767718080682e+17, 1.27767718090682e+17, 1.27767718100682e+17, 1.277677181092758e+17, 1.277677181183383e+17, 1.27767718130682e+17, 1.27767718140682e+17, 1.277677181494321e+17, 1.27767718160682e+17, 1.27767718168182e+17, 1.27767718180682e+17, 1.277677181872445e+17, 1.27767718200682e+17, 1.27767718210682e+17, 1.277677182192758e+17, 1.277677182306821e+17, 1.277677182374008e+17, 1.277677182464634e+17, 1.27767718260682e+17, 1.27767718270682e+17, 1.277677182794319e+17, 1.27767718290682e+17, 1.277677182974007e+17, 1.277677183066195e+17, 1.27767718320682e+17, 1.27767718330682e+17, 1.277677183394321e+17},
			             {1.27767691700682e+17, 1.27767691710682e+17, 1.27767691720682e+17, 1.27767691730682e+17, 1.27767691740682e+17, 1.277676917506821e+17, 1.27767691760682e+17, 1.27767691770682e+17, 1.27767691780682e+17, 1.27767691790682e+17, 1.27767691800682e+17, 1.27767691810682e+17, 1.27767691820682e+17, 1.27767691830682e+17, 1.27767691840682e+17, 1.27767691850682e+17, 1.27767691860682e+17, 1.27767691870682e+17, 1.27767691880682e+17, 1.27767691890682e+17, 1.27767691900682e+17, 1.27767691910682e+17, 1.27767691920682e+17, 1.27767691930682e+17, 1.27767691940682e+17, 1.27767691950682e+17, 1.27767691960682e+17, 1.27767691970682e+17, 1.27767691980682e+17, 1.27767691990682e+17, 1.27767692000682e+17, 1.27767692010682e+17, 1.27767692020682e+17, 1.27767692030682e+17, 1.27767692040682e+17, 1.27767692050682e+17, 1.27767692060682e+17, 1.27767692070682e+17, 1.27767692080682e+17, 1.27767692090682e+17, 1.27767692100682e+17, 1.27767692110682e+17, 1.277676921206821e+17, 1.27767692130682e+17, 1.27767692140682e+17, 1.27767692150682e+17, 1.27767692160682e+17, 1.27767692170682e+17},
			             {1.27767692400682e+17, 1.27767692410682e+17, 1.27767692420682e+17, 1.27767692430682e+17, 1.27767692440682e+17, 1.27767692450682e+17, 1.27767692460682e+17, 1.27767692470682e+17, 1.27767692480682e+17, 1.27767692490682e+17, 1.27767692500682e+17, 1.27767692510682e+17, 1.27767692520682e+17, 1.27767692530682e+17, 1.27767692540682e+17, 1.27767692550682e+17, 1.27767692560682e+17, 1.27767692570682e+17, 1.27767692580682e+17, 1.27767692590682e+17, 1.27767692600682e+17, 1.27767692610682e+17},
			             {1.27767693370682e+17, 1.27767693380682e+17, 1.27767693390682e+17, 1.27767693400682e+17, 1.27767693410682e+17, 1.27767693420682e+17, 1.27767693430682e+17, 1.27767693440682e+17, 1.27767693450682e+17, 1.27767693460682e+17, 1.27767693470682e+17, 1.27767693480682e+17, 1.27767693490682e+17, 1.27767693500682e+17, 1.27767693510682e+17, 1.27767693520682e+17, 1.277676935306821e+17, 1.27767693540682e+17, 1.27767693550682e+17, 1.27767693560682e+17, 1.27767693570682e+17, 1.27767693580682e+17, 1.27767693590682e+17, 1.27767693600682e+17, 1.27767693610682e+17, 1.27767693620682e+17, 1.27767693630682e+17},
			             {1.27767691610682e+17, 1.27767691620682e+17, 1.27767691630682e+17, 1.27767691640682e+17, 1.27767691650682e+17, 1.27767691660682e+17, 1.27767691670682e+17, 1.27767691680682e+17, 1.27767691690682e+17, 1.27767691700682e+17, 1.27767691710682e+17, 1.27767691720682e+17, 1.27767691730682e+17, 1.27767691740682e+17, 1.277676917506821e+17, 1.27767691760682e+17, 1.27767691770682e+17, 1.27767691780682e+17, 1.27767691790682e+17, 1.27767691800682e+17, 1.27767691810682e+17, 1.27767691820682e+17, 1.27767691830682e+17, 1.27767691840682e+17, 1.27767691850682e+17, 1.27767691860682e+17, 1.27767691870682e+17, 1.27767691880682e+17, 1.27767691890682e+17, 1.27767691900682e+17, 1.27767691910682e+17, 1.27767691920682e+17, 1.27767691930682e+17, 1.27767691940682e+17, 1.27767691950682e+17, 1.27767691960682e+17, 1.27767691970682e+17, 1.27767691980682e+17, 1.27767691990682e+17, 1.27767692000682e+17, 1.27767692010682e+17, 1.27767692020682e+17, 1.27767692030682e+17, 1.27767692040682e+17, 1.27767692050682e+17, 1.27767692060682e+17, 1.27767692070682e+17, 1.27767692080682e+17, 1.27767692090682e+17, 1.27767692100682e+17, 1.27767692110682e+17, 1.277676921206821e+17, 1.27767692130682e+17, 1.27767692140682e+17, 1.27767692150682e+17, 1.27767692160682e+17, 1.27767692170682e+17, 1.27767692180682e+17, 1.27767692190682e+17, 1.27767692200682e+17, 1.27767692210682e+17, 1.27767692220682e+17, 1.27767692230682e+17, 1.27767692240682e+17, 1.27767692250682e+17, 1.27767692260682e+17, 1.27767692270682e+17, 1.27767692280682e+17, 1.27767692290682e+17, 1.27767692300682e+17, 1.27767692310682e+17, 1.27767692320682e+17, 1.27767692330682e+17, 1.27767692340682e+17, 1.27767692350682e+17, 1.27767692360682e+17, 1.27767692370682e+17},
			             {1.27767688240682e+17, 1.27767688250682e+17, 1.27767688260682e+17, 1.27767688270682e+17, 1.27767688280682e+17, 1.27767688290682e+17, 1.277676883006821e+17, 1.27767688310682e+17, 1.27767688320682e+17, 1.27767688330682e+17, 1.27767688340682e+17, 1.27767688350682e+17, 1.27767688360682e+17, 1.27767688370682e+17, 1.27767688380682e+17, 1.27767688390682e+17, 1.27767688400682e+17, 1.27767688410682e+17, 1.27767688420682e+17, 1.27767688430682e+17, 1.27767688440682e+17, 1.27767688450682e+17, 1.27767688460682e+17, 1.27767688470682e+17, 1.27767688480682e+17, 1.27767688490682e+17, 1.27767688500682e+17, 1.27767688510682e+17, 1.27767688520682e+17, 1.27767688530682e+17, 1.27767688540682e+17, 1.27767688550682e+17, 1.277676885606821e+17, 1.27767688570682e+17, 1.27767688580682e+17, 1.27767688590682e+17, 1.27767688600682e+17, 1.27767688610682e+17, 1.27767688620682e+17, 1.27767688630682e+17, 1.27767688640682e+17, 1.27767688650682e+17, 1.27767688660682e+17, 1.27767688670682e+17, 1.27767688680682e+17, 1.27767688690682e+17, 1.27767688700682e+17, 1.27767688710682e+17, 1.27767688720682e+17, 1.27767688730682e+17, 1.27767688740682e+17, 1.27767688750682e+17, 1.27767688760682e+17, 1.27767688770682e+17, 1.27767688780682e+17, 1.27767688790682e+17, 1.27767688800682e+17, 1.27767688810682e+17, 1.277676888206821e+17, 1.27767688830682e+17, 1.27767688840682e+17, 1.27767688850682e+17, 1.27767688860682e+17, 1.27767688870682e+17, 1.27767688880682e+17, 1.27767688890682e+17, 1.27767688900682e+17, 1.27767688910682e+17, 1.27767688920682e+17, 1.27767688930682e+17, 1.27767688940682e+17, 1.27767688950682e+17, 1.27767688960682e+17, 1.27767688970682e+17, 1.27767688980682e+17, 1.27767688990682e+17, 1.27767689000682e+17, 1.27767689010682e+17, 1.27767689020682e+17, 1.27767689030682e+17, 1.27767689040682e+17, 1.27767689050682e+17, 1.27767689060682e+17, 1.27767689070682e+17, 1.27767689080682e+17, 1.27767689090682e+17, 1.27767689100682e+17, 1.27767689110682e+17, 1.27767689120682e+17, 1.27767689130682e+17, 1.27767689140682e+17, 1.27767689150682e+17, 1.27767689160682e+17, 1.27767689170682e+17, 1.27767689180682e+17, 1.277676891906821e+17, 1.27767689200682e+17, 1.27767689210682e+17, 1.27767689220682e+17, 1.27767689230682e+17, 1.27767689240682e+17, 1.27767689250682e+17, 1.27767689260682e+17, 1.27767689270682e+17, 1.27767689280682e+17, 1.27767689290682e+17, 1.27767689300682e+17, 1.27767689310682e+17, 1.27767689320682e+17, 1.27767689330682e+17, 1.27767689340682e+17, 1.27767689350682e+17, 1.27767689360682e+17, 1.27767689370682e+17, 1.27767689380682e+17, 1.27767689390682e+17, 1.27767689400682e+17, 1.27767689410682e+17, 1.27767689420682e+17, 1.27767689430682e+17, 1.27767689440682e+17, 1.277676894506821e+17, 1.27767689460682e+17, 1.27767689470682e+17, 1.27767689480682e+17, 1.27767689490682e+17, 1.27767689500682e+17, 1.27767689510682e+17, 1.27767689520682e+17, 1.27767689530682e+17, 1.27767689540682e+17, 1.27767689550682e+17, 1.27767689560682e+17, 1.27767689570682e+17, 1.27767689580682e+17, 1.27767689590682e+17, 1.27767689600682e+17, 1.27767689610682e+17, 1.27767689620682e+17, 1.27767689630682e+17, 1.27767689640682e+17, 1.27767689650682e+17, 1.27767689660682e+17, 1.27767689670682e+17, 1.27767689680682e+17, 1.27767689690682e+17, 1.27767689700682e+17, 1.277676897106821e+17, 1.27767689720682e+17, 1.27767689730682e+17, 1.27767689740682e+17, 1.27767689750682e+17, 1.27767689760682e+17, 1.27767689770682e+17, 1.27767689780682e+17, 1.27767689790682e+17, 1.27767689800682e+17, 1.27767689810682e+17, 1.27767689820682e+17, 1.27767689830682e+17, 1.27767689840682e+17, 1.27767689850682e+17, 1.27767689860682e+17, 1.27767689870682e+17, 1.27767689880682e+17, 1.27767689890682e+17, 1.27767689900682e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}};
		}
	}
}
