netcdf mask {
	:date_created = "20200811T114628";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200811T114628";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 11;
			channels = 6;
			categories = 35;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  172.4, 181.1, 178.8, 186.6, 179.3, 130.3, 120.1, 112.4, 107.0, 102.6,  99.1;
			max_depth =  197.8, 189.2, 185.6, 198.6, 185.7, 205.7, 152.7, 144.6, 166.3, 153.0, 146.4;
			start_time = 127767706080681984, 127767702330681984, 127767702600681984, 127767703200681984, 127767703100681984, 127767707040681984, 127767691700681984, 127767692400681984, 127767693370681984, 127767691610681984, 127767688240681984;
			end_time = 127767706210681984, 127767702430681984, 127767702640681984, 127767703240681984, 127767703160681984, 127767718339432064, 127767692170681984, 127767692610681984, 127767693630681984, 127767692370681984, 127767689900681984;
			region_id = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11;
			region_name = "Layer1","Layer2","Layer3","Layer4","Layer5","Layer6","Layer7","Layer8","Layer9","Layer10","Layer11";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "", "", "", "", "", "", "", "";
			region_category_names = "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "21", "12", "12", "12", "12", "12", "12", "12", "12", "12", "12", "12", "12";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35;
			region_type = analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis, analysis;
			channel_names = "18", "38", "70", "120", "200", "364";
			region_channels = 0, 16, 16, 16, 16, 16, 63, 63, 63, 63, 63;
			mask_times = {1.27767706080682e+17, 1.27767706090682e+17, 1.27767706100682e+17, 1.27767706110682e+17, 1.27767706120682e+17, 1.27767706130682e+17, 1.277677061406821e+17, 1.27767706150682e+17, 1.27767706160682e+17, 1.27767706170682e+17, 1.27767706180682e+17, 1.27767706190682e+17, 1.27767706200682e+17, 1.27767706210682e+17},
			             {1.27767702330682e+17, 1.27767702340682e+17, 1.27767702350682e+17, 1.27767702360682e+17, 1.27767702370682e+17, 1.27767702380682e+17, 1.27767702390682e+17, 1.27767702400682e+17, 1.27767702410682e+17, 1.27767702420682e+17, 1.27767702430682e+17},
			             {1.27767702600682e+17, 1.27767702610682e+17, 1.27767702620682e+17, 1.27767702630682e+17, 1.27767702640682e+17},
			             {1.27767703200682e+17, 1.277677032106821e+17, 1.27767703220682e+17, 1.27767703230682e+17, 1.27767703240682e+17},
			             {1.27767703100682e+17, 1.27767703110682e+17, 1.27767703120682e+17, 1.27767703130682e+17, 1.27767703140682e+17, 1.27767703150682e+17, 1.27767703160682e+17},
			             {1.27767707040682e+17, 1.27767707050682e+17, 1.27767707060682e+17, 1.27767707070682e+17, 1.27767707080682e+17, 1.27767707090682e+17, 1.27767707100682e+17, 1.27767707110682e+17, 1.27767707120682e+17, 1.27767707130682e+17, 1.27767707140682e+17, 1.27767707150682e+17, 1.27767707160682e+17, 1.27767707170682e+17, 1.27767707180682e+17, 1.27767707190682e+17, 1.27767707200682e+17, 1.27767707210682e+17, 1.27767707220682e+17, 1.27767707230682e+17, 1.27767707240682e+17, 1.27767707250682e+17, 1.27767707260682e+17, 1.27767707270682e+17, 1.27767707280682e+17, 1.27767707290682e+17, 1.27767707300682e+17, 1.27767707310682e+17, 1.27767707320682e+17, 1.27767707330682e+17, 1.27767707340682e+17, 1.27767707350682e+17, 1.27767707360682e+17, 1.27767707370682e+17, 1.27767707380682e+17, 1.27767707390682e+17, 1.27767707400682e+17, 1.27767707410682e+17, 1.27767707420682e+17, 1.27767707430682e+17, 1.27767707440682e+17, 1.27767707450682e+17, 1.27767707460682e+17, 1.27767707470682e+17, 1.27767707480682e+17, 1.27767707490682e+17, 1.27767707500682e+17, 1.27767707510682e+17, 1.27767707520682e+17, 1.27767707530682e+17, 1.27767707540682e+17, 1.27767707550682e+17, 1.27767707560682e+17, 1.27767707570682e+17, 1.27767707580682e+17, 1.27767707590682e+17, 1.27767707600682e+17, 1.27767707610682e+17, 1.27767707620682e+17, 1.27767707630682e+17, 1.27767707640682e+17, 1.27767707650682e+17, 1.277677076606821e+17, 1.27767707670682e+17, 1.27767707680682e+17, 1.27767707690682e+17, 1.27767707700682e+17, 1.27767707710682e+17, 1.27767707720682e+17, 1.27767707730682e+17, 1.27767707740682e+17, 1.27767707750682e+17, 1.27767707760682e+17, 1.27767707770682e+17, 1.27767707780682e+17, 1.27767707790682e+17, 1.27767707800682e+17, 1.27767707810682e+17, 1.27767707820682e+17, 1.27767707830682e+17, 1.27767707840682e+17, 1.27767707850682e+17, 1.27767707860682e+17, 1.27767707870682e+17, 1.27767707880682e+17, 1.27767707890682e+17, 1.27767707900682e+17, 1.27767707910682e+17, 1.277677079206821e+17, 1.27767707930682e+17, 1.27767707940682e+17, 1.27767707950682e+17, 1.27767707960682e+17, 1.27767707970682e+17, 1.27767707980682e+17, 1.27767707990682e+17, 1.27767708000682e+17, 1.27767708010682e+17, 1.27767708020682e+17, 1.27767708030682e+17, 1.27767708040682e+17, 1.27767708050682e+17, 1.27767708060682e+17, 1.27767708070682e+17, 1.27767708080682e+17, 1.27767708090682e+17, 1.27767708100682e+17, 1.27767708110682e+17, 1.27767708120682e+17, 1.27767708130682e+17, 1.27767708140682e+17, 1.27767708150682e+17, 1.27767708160682e+17, 1.27767708170682e+17, 1.277677081806821e+17, 1.27767708190682e+17, 1.27767708200682e+17, 1.27767708210682e+17, 1.27767708220682e+17, 1.27767708230682e+17, 1.27767708240682e+17, 1.27767708250682e+17, 1.27767708260682e+17, 1.27767708270682e+17, 1.27767708280682e+17, 1.27767708290682e+17, 1.27767708300682e+17, 1.27767708310682e+17, 1.27767708320682e+17, 1.27767708330682e+17, 1.27767708340682e+17, 1.27767708350682e+17, 1.27767708360682e+17, 1.27767708370682e+17, 1.27767708380682e+17, 1.27767708390682e+17, 1.27767708400682e+17, 1.27767708410682e+17, 1.27767708420682e+17, 1.27767708430682e+17, 1.27767708440682e+17, 1.27767708450682e+17, 1.27767708460682e+17, 1.27767708470682e+17, 1.27767708480682e+17, 1.27767708490682e+17, 1.27767708500682e+17, 1.27767708510682e+17, 1.27767708520682e+17, 1.27767708530682e+17, 1.27767708540682e+17, 1.277677085506821e+17, 1.27767708560682e+17, 1.27767708570682e+17, 1.27767708580682e+17, 1.27767708590682e+17, 1.27767708600682e+17, 1.27767708610682e+17, 1.27767708620682e+17, 1.27767708630682e+17, 1.27767708640682e+17, 1.27767708650682e+17, 1.27767708660682e+17, 1.27767708670682e+17, 1.27767708680682e+17, 1.27767708690682e+17, 1.27767708700682e+17, 1.27767708710682e+17, 1.27767708720682e+17, 1.27767708730682e+17, 1.27767708740682e+17, 1.27767708750682e+17, 1.27767708760682e+17, 1.27767708770682e+17, 1.27767708780682e+17, 1.27767708790682e+17, 1.27767708800682e+17, 1.277677088106821e+17, 1.27767708820682e+17, 1.27767708830682e+17, 1.27767708840682e+17, 1.27767708850682e+17, 1.27767708860682e+17, 1.27767708870682e+17, 1.27767708880682e+17, 1.27767708890682e+17, 1.27767708900682e+17, 1.27767708910682e+17, 1.27767708920682e+17, 1.27767708930682e+17, 1.27767708940682e+17, 1.27767708950682e+17, 1.27767708960682e+17, 1.27767708970682e+17, 1.27767708980682e+17, 1.27767708990682e+17, 1.27767709000682e+17, 1.27767709010682e+17, 1.27767709020682e+17, 1.27767709030682e+17, 1.27767709040682e+17, 1.27767709050682e+17, 1.27767709060682e+17, 1.277677090706821e+17, 1.27767709080682e+17, 1.27767709090682e+17, 1.27767709100682e+17, 1.27767709110682e+17, 1.27767709120682e+17, 1.27767709130682e+17, 1.27767709140682e+17, 1.27767709150682e+17, 1.27767709160682e+17, 1.27767709170682e+17, 1.27767709180682e+17, 1.27767709190682e+17, 1.27767709200682e+17, 1.27767709210682e+17, 1.27767709220682e+17, 1.27767709230682e+17, 1.27767709240682e+17, 1.27767709250682e+17, 1.27767709260682e+17, 1.27767709270682e+17, 1.27767709280682e+17, 1.27767709290682e+17, 1.27767709300682e+17, 1.27767709310682e+17, 1.27767709320682e+17, 1.27767709330682e+17, 1.27767709340682e+17, 1.27767709350682e+17, 1.27767709360682e+17, 1.27767709370682e+17, 1.27767709380682e+17, 1.27767709390682e+17, 1.27767709420682e+17, 1.27767709430682e+17, 1.277677094406821e+17, 1.27767709450682e+17, 1.27767709460682e+17, 1.27767709470682e+17, 1.27767709480682e+17, 1.27767709490682e+17, 1.27767709500682e+17, 1.27767709510682e+17, 1.27767709520682e+17, 1.27767709530682e+17, 1.27767709540682e+17, 1.27767709550682e+17, 1.27767709560682e+17, 1.27767709570682e+17, 1.27767709580682e+17, 1.27767709590682e+17, 1.27767709600682e+17, 1.27767709610682e+17, 1.27767709620682e+17, 1.27767709630682e+17, 1.27767709640682e+17, 1.27767709650682e+17, 1.27767709660682e+17, 1.27767709670682e+17, 1.27767709680682e+17, 1.27767709690682e+17, 1.277677097006821e+17, 1.27767709710682e+17, 1.27767709720682e+17, 1.27767709730682e+17, 1.27767709740682e+17, 1.27767709750682e+17, 1.27767709760682e+17, 1.27767709770682e+17, 1.27767709780682e+17, 1.27767709790682e+17, 1.27767709800682e+17, 1.27767709810682e+17, 1.27767709820682e+17, 1.27767709830682e+17, 1.27767709840682e+17, 1.27767709850682e+17, 1.27767709860682e+17, 1.27767709870682e+17, 1.27767709880682e+17, 1.27767709890682e+17, 1.27767709900682e+17, 1.27767709910682e+17, 1.27767709920682e+17, 1.27767709930682e+17, 1.27767709940682e+17, 1.27767709950682e+17, 1.277677099606821e+17, 1.27767709970682e+17, 1.27767709980682e+17, 1.27767709990682e+17, 1.27767710000682e+17, 1.27767710010682e+17, 1.27767710020682e+17, 1.27767710030682e+17, 1.27767710040682e+17, 1.27767710050682e+17, 1.27767710060682e+17, 1.27767710070682e+17, 1.27767710080682e+17, 1.27767710090682e+17, 1.27767710100682e+17, 1.27767710110682e+17, 1.27767710120682e+17, 1.27767710130682e+17, 1.27767710140682e+17, 1.27767710150682e+17, 1.27767710160682e+17, 1.27767710170682e+17, 1.27767710180682e+17, 1.27767710190682e+17, 1.27767710200682e+17, 1.27767710210682e+17, 1.27767710220682e+17, 1.27767710230682e+17, 1.27767710240682e+17, 1.27767710250682e+17, 1.27767710260682e+17, 1.27767710270682e+17, 1.27767710280682e+17, 1.27767710290682e+17, 1.27767710300682e+17, 1.27767710310682e+17, 1.27767710320682e+17, 1.277677103306821e+17, 1.27767710340682e+17, 1.27767710350682e+17, 1.27767710360682e+17, 1.27767710370682e+17, 1.27767710380682e+17, 1.27767710390682e+17, 1.27767710400682e+17, 1.27767710410682e+17, 1.27767710420682e+17, 1.27767710430682e+17, 1.27767710440682e+17, 1.27767710450682e+17, 1.27767710460682e+17, 1.27767710470682e+17, 1.27767710480682e+17, 1.27767710490682e+17, 1.27767710500682e+17, 1.27767710510682e+17, 1.27767710520682e+17, 1.27767710530682e+17, 1.27767710540682e+17, 1.27767710550682e+17, 1.27767710560682e+17, 1.27767710570682e+17, 1.27767710580682e+17, 1.277677105906821e+17, 1.27767710600682e+17, 1.27767710610682e+17, 1.27767710620682e+17, 1.27767710630682e+17, 1.27767710640682e+17, 1.27767710650682e+17, 1.27767710660682e+17, 1.27767710670682e+17, 1.27767710680682e+17, 1.27767710690682e+17, 1.27767710700682e+17, 1.27767710710682e+17, 1.27767710720682e+17, 1.27767710730682e+17, 1.27767710740682e+17, 1.27767710750682e+17, 1.27767710760682e+17, 1.27767710770682e+17, 1.27767710780682e+17, 1.27767710790682e+17, 1.27767710800682e+17, 1.27767710810682e+17, 1.27767710820682e+17, 1.27767710830682e+17, 1.27767710840682e+17, 1.277677108506821e+17, 1.27767710860682e+17, 1.277677108678696e+17, 1.27767710880682e+17, 1.277677108903695e+17, 1.277677108975571e+17, 1.27767710910682e+17, 1.27767710920682e+17, 1.277677109297445e+17, 1.277677109359945e+17, 1.27767710950682e+17, 1.27767710960682e+17, 1.27767710970682e+17, 1.27767710980682e+17, 1.27767710990682e+17, 1.27767711000682e+17, 1.277677110070883e+17, 1.277677110167757e+17, 1.27767711030682e+17, 1.27767711040682e+17, 1.27767711050682e+17, 1.27767711060682e+17, 1.277677110699008e+17, 1.27767711080682e+17, 1.27767711090682e+17, 1.27767711100682e+17, 1.27767711110682e+17, 1.277677111202132e+17, 1.27767711130682e+17, 1.27767711140682e+17, 1.27767711150682e+17, 1.27767711160682e+17, 1.27767711170057e+17, 1.27767711180682e+17, 1.27767711190682e+17, 1.27767711200682e+17, 1.27767711210682e+17, 1.277677112202132e+17, 1.27767711230682e+17, 1.27767711240682e+17, 1.27767711250682e+17, 1.27767711260682e+17, 1.277677112694319e+17, 1.27767711280682e+17, 1.27767711290682e+17, 1.27767711300682e+17, 1.27767711310682e+17, 1.277677113195882e+17, 1.27767711330682e+17, 1.27767711340682e+17, 1.27767711350682e+17, 1.27767711360682e+17, 1.27767711370682e+17, 1.277677113803695e+17, 1.27767711390682e+17, 1.27767711400682e+17, 1.27767711410682e+17, 1.27767711420682e+17, 1.277677114295882e+17, 1.27767711440682e+17, 1.27767711450682e+17, 1.27767711460682e+17, 1.27767711470682e+17, 1.277677114792756e+17, 1.27767711490682e+17, 1.27767711500682e+17, 1.27767711510682e+17, 1.27767711520682e+17, 1.277677115295882e+17, 1.27767711540682e+17, 1.27767711550682e+17, 1.27767711560682e+17, 1.27767711570682e+17, 1.277677115797445e+17, 1.27767711590682e+17, 1.27767711600682e+17, 1.27767711610682e+17, 1.27767711620682e+17, 1.277677116295884e+17, 1.27767711640682e+17, 1.27767711650682e+17, 1.27767711660682e+17, 1.27767711670682e+17, 1.277677116799008e+17, 1.27767711690682e+17, 1.27767711700682e+17, 1.27767711710682e+17, 1.27767711720682e+17, 1.27767711730057e+17, 1.277677117406821e+17, 1.27767711750682e+17, 1.27767711760682e+17, 1.27767711770682e+17, 1.277677117799007e+17, 1.27767711790682e+17, 1.27767711800682e+17, 1.27767711810682e+17, 1.27767711820682e+17, 1.277677118302132e+17, 1.27767711840682e+17, 1.27767711850682e+17, 1.27767711860682e+17, 1.27767711870682e+17, 1.277677118792758e+17, 1.27767711890682e+17, 1.27767711900682e+17, 1.27767711910682e+17, 1.27767711920682e+17, 1.27767711930682e+17, 1.27767711940682e+17, 1.27767711950682e+17, 1.27767711960682e+17, 1.27767711970682e+17, 1.277677119803695e+17, 1.277677119903695e+17, 1.277677120006821e+17, 1.27767712010682e+17, 1.27767712020682e+17, 1.27767712030682e+17, 1.277677120395884e+17, 1.27767712050682e+17, 1.27767712060682e+17, 1.27767712070682e+17, 1.27767712080682e+17, 1.277677120902132e+17, 1.27767712100682e+17, 1.27767712110682e+17, 1.27767712120682e+17, 1.27767712130682e+17, 1.277677121402132e+17, 1.27767712150682e+17, 1.27767712160682e+17, 1.27767712170682e+17, 1.27767712180682e+17, 1.277677121895882e+17, 1.27767712200682e+17, 1.27767712210682e+17, 1.27767712220682e+17, 1.27767712230682e+17, 1.277677122397445e+17, 1.27767712250682e+17, 1.27767712260682e+17, 1.27767712270682e+17, 1.27767712280682e+17, 1.277677122899008e+17, 1.27767712300682e+17, 1.27767712310682e+17, 1.27767712320682e+17, 1.27767712330682e+17, 1.277677123397445e+17, 1.27767712350682e+17, 1.27767712360682e+17, 1.277677123706821e+17, 1.27767712380682e+17, 1.27767712390057e+17, 1.27767712400682e+17, 1.27767712410682e+17, 1.27767712420682e+17, 1.27767712430682e+17, 1.277677124397444e+17, 1.27767712450682e+17, 1.27767712460682e+17, 1.27767712470682e+17, 1.277677124799007e+17, 1.27767712490682e+17, 1.27767712500682e+17, 1.27767712510682e+17, 1.27767712520057e+17, 1.27767712530682e+17, 1.27767712540682e+17, 1.27767712550682e+17, 1.27767712560057e+17, 1.27767712570682e+17, 1.27767712580682e+17, 1.27767712590682e+17, 1.277677126002132e+17, 1.27767712610682e+17, 1.27767712620682e+17, 1.277677126306821e+17, 1.277677126394319e+17, 1.27767712650682e+17, 1.27767712660682e+17, 1.27767712670682e+17, 1.277677126794319e+17, 1.27767712690682e+17, 1.27767712700682e+17, 1.27767712710682e+17, 1.277677127202132e+17, 1.27767712730682e+17, 1.27767712740682e+17, 1.27767712750682e+17, 1.277677127594321e+17, 1.27767712770682e+17, 1.27767712780682e+17, 1.27767712790682e+17, 1.277677127995884e+17, 1.27767712810682e+17, 1.27767712820682e+17, 1.27767712830682e+17, 1.277677128397445e+17, 1.27767712850682e+17, 1.27767712860682e+17, 1.27767712870682e+17, 1.277677128795882e+17, 1.277677128906821e+17, 1.27767712900682e+17, 1.27767712910682e+17, 1.277677129195882e+17, 1.27767712930682e+17, 1.27767712940682e+17, 1.27767712950682e+17, 1.277677129597444e+17, 1.27767712970682e+17, 1.27767712980682e+17, 1.27767712990682e+17, 1.277677129999007e+17, 1.27767713010682e+17, 1.27767713020682e+17, 1.27767713030682e+17, 1.277677130397445e+17, 1.27767713050682e+17, 1.27767713060682e+17, 1.27767713070682e+17, 1.277677130799008e+17, 1.27767713090682e+17, 1.27767713100682e+17, 1.27767713110682e+17, 1.277677131199008e+17, 1.27767713130682e+17, 1.27767713140682e+17, 1.27767713150682e+17, 1.27767713160057e+17, 1.27767713170682e+17, 1.27767713180682e+17, 1.27767713190682e+17, 1.277677131992758e+17, 1.27767713210682e+17, 1.27767713220682e+17, 1.27767713230682e+17, 1.277677132400571e+17, 1.27767713250682e+17, 1.277677132606821e+17, 1.27767713270682e+17, 1.277677132802132e+17, 1.27767713290682e+17, 1.27767713300682e+17, 1.27767713310682e+17, 1.277677133192758e+17, 1.27767713330682e+17, 1.27767713340682e+17, 1.27767713350682e+17, 1.277677133595882e+17, 1.27767713370682e+17, 1.27767713380682e+17, 1.27767713390682e+17, 1.277677133994319e+17, 1.27767713410682e+17, 1.27767713420682e+17, 1.27767713430682e+17, 1.277677134394321e+17, 1.27767713450682e+17, 1.27767713460682e+17, 1.27767713470682e+17, 1.277677134795882e+17, 1.27767713490682e+17, 1.27767713500682e+17, 1.27767713510682e+17, 1.277677135202132e+17, 1.27767713530682e+17, 1.27767713540682e+17, 1.27767713550682e+17, 1.277677135595884e+17, 1.27767713570682e+17, 1.27767713580682e+17, 1.27767713590682e+17, 1.277677135995882e+17, 1.27767713610682e+17, 1.27767713620682e+17, 1.27767713630682e+17, 1.277677136397445e+17, 1.27767713650682e+17, 1.27767713660682e+17, 1.27767713670682e+17, 1.277677136799008e+17, 1.27767713690682e+17, 1.27767713700682e+17, 1.27767713710682e+17, 1.277677137197445e+17, 1.27767713730682e+17, 1.27767713740682e+17, 1.27767713750682e+17, 1.277677137599007e+17, 1.27767713770682e+17, 1.277677137806821e+17, 1.27767713790682e+17, 1.27767713800057e+17, 1.27767713810682e+17, 1.27767713820682e+17, 1.27767713830682e+17, 1.277677138402132e+17, 1.27767713850682e+17, 1.27767713860682e+17, 1.27767713870682e+17, 1.27767713880057e+17, 1.27767713890682e+17, 1.27767713900682e+17, 1.27767713910682e+17, 1.277677139202132e+17, 1.27767713930682e+17, 1.27767713940682e+17, 1.27767713950682e+17, 1.277677139592758e+17, 1.27767713970682e+17, 1.27767713980682e+17, 1.27767713990682e+17, 1.277677139994321e+17, 1.27767714010682e+17, 1.27767714020682e+17, 1.27767714030682e+17, 1.277677140402132e+17, 1.27767714050682e+17, 1.27767714060682e+17, 1.27767714070682e+17, 1.277677140794319e+17, 1.27767714090682e+17, 1.27767714100682e+17, 1.27767714110682e+17, 1.27767714120057e+17, 1.27767714130682e+17, 1.27767714140682e+17, 1.27767714150682e+17, 1.277677141602132e+17, 1.27767714170682e+17, 1.27767714180682e+17, 1.27767714190682e+17, 1.277677141994319e+17, 1.27767714210682e+17, 1.27767714220682e+17, 1.27767714230682e+17, 1.277677142395882e+17, 1.27767714250682e+17, 1.27767714260682e+17, 1.27767714270682e+17, 1.277677142797445e+17, 1.27767714290682e+17, 1.27767714300682e+17, 1.27767714310682e+17, 1.277677143199008e+17, 1.27767714330682e+17, 1.27767714340682e+17, 1.27767714350682e+17, 1.277677143594319e+17, 1.27767714370682e+17, 1.27767714380682e+17, 1.27767714390682e+17, 1.277677143997445e+17, 1.277677144106821e+17, 1.27767714420682e+17, 1.27767714430682e+17, 1.277677144399008e+17, 1.27767714450682e+17, 1.27767714460682e+17, 1.27767714470682e+17, 1.277677144800571e+17, 1.27767714490682e+17, 1.27767714500682e+17, 1.27767714510682e+17, 1.277677145194321e+17, 1.27767714530682e+17, 1.27767714540682e+17, 1.27767714550682e+17, 1.27767714560057e+17, 1.27767714570682e+17, 1.27767714580682e+17, 1.27767714590682e+17, 1.277677146002132e+17, 1.27767714610682e+17, 1.27767714620682e+17, 1.27767714630682e+17, 1.277677146392758e+17, 1.27767714650682e+17, 1.27767714660682e+17, 1.277677146706821e+17, 1.277677146794319e+17, 1.27767714690682e+17, 1.27767714700682e+17, 1.27767714710682e+17, 1.277677147202132e+17, 1.27767714730682e+17, 1.27767714740682e+17, 1.27767714750682e+17, 1.277677147592758e+17, 1.27767714770682e+17, 1.27767714780682e+17, 1.27767714790682e+17, 1.277677147994321e+17, 1.27767714810682e+17, 1.27767714820682e+17, 1.27767714830682e+17, 1.277677148395884e+17, 1.27767714850682e+17, 1.27767714860682e+17, 1.27767714870682e+17, 1.277677148794319e+17, 1.27767714890682e+17, 1.27767714900682e+17, 1.27767714910682e+17, 1.277677149195882e+17, 1.277677149306821e+17, 1.27767714940682e+17, 1.277677149486508e+17, 1.277677149586508e+17, 1.27767714970682e+17, 1.27767714980682e+17, 1.27767714990682e+17, 1.277677149999008e+17, 1.27767715010682e+17, 1.27767715020682e+17, 1.27767715030682e+17, 1.277677150395884e+17, 1.27767715050682e+17, 1.27767715060682e+17, 1.27767715070682e+17, 1.277677150797445e+17, 1.27767715090682e+17, 1.27767715100682e+17, 1.27767715110682e+17, 1.277677151199008e+17, 1.27767715130682e+17, 1.27767715140682e+17, 1.27767715150682e+17, 1.27767715160057e+17, 1.27767715170682e+17, 1.27767715180682e+17, 1.27767715190682e+17, 1.277677151999008e+17, 1.27767715210682e+17, 1.27767715220682e+17, 1.27767715230682e+17, 1.277677152399008e+17, 1.27767715250682e+17, 1.27767715260682e+17, 1.27767715270682e+17, 1.277677152799007e+17, 1.27767715290682e+17, 1.277677153006821e+17, 1.27767715310682e+17, 1.27767715320057e+17, 1.27767715330682e+17, 1.27767715340682e+17, 1.27767715350682e+17, 1.277677153602132e+17, 1.27767715370682e+17, 1.27767715380682e+17, 1.27767715390682e+17, 1.277677153992758e+17, 1.27767715410682e+17, 1.27767715420682e+17, 1.27767715430682e+17, 1.277677154394319e+17, 1.27767715450682e+17, 1.27767715460682e+17, 1.27767715470682e+17, 1.277677154800571e+17, 1.27767715490682e+17, 1.27767715500682e+17, 1.27767715510682e+17, 1.277677155194321e+17, 1.27767715530682e+17, 1.27767715540682e+17, 1.27767715550682e+17, 1.277677155595884e+17, 1.27767715570682e+17, 1.27767715580682e+17, 1.27767715590682e+17, 1.277677155997445e+17, 1.27767715610682e+17, 1.27767715620682e+17, 1.27767715630682e+17, 1.277677156397445e+17, 1.27767715650682e+17, 1.27767715660682e+17, 1.27767715670682e+17, 1.277677156795882e+17, 1.27767715690682e+17, 1.27767715700682e+17, 1.27767715710682e+17, 1.277677157197445e+17, 1.27767715730682e+17, 1.27767715740682e+17, 1.27767715750682e+17, 1.277677157599008e+17, 1.27767715770682e+17, 1.27767715780682e+17, 1.27767715790682e+17, 1.27767715800682e+17, 1.27767715810682e+17, 1.277677158206821e+17, 1.27767715830682e+17, 1.277677158399008e+17, 1.27767715850682e+17, 1.27767715860682e+17, 1.27767715870682e+17, 1.27767715880057e+17, 1.27767715890682e+17, 1.27767715900682e+17, 1.27767715910682e+17, 1.277677159202132e+17, 1.27767715930682e+17, 1.27767715940682e+17, 1.27767715950682e+17, 1.277677159597445e+17, 1.27767715970682e+17, 1.27767715980682e+17, 1.27767715990682e+17, 1.277677160000571e+17, 1.27767716010682e+17, 1.27767716020682e+17, 1.27767716030682e+17, 1.277677160402132e+17, 1.27767716050682e+17, 1.27767716060682e+17, 1.27767716070682e+17, 1.277677160794321e+17, 1.27767716090682e+17, 1.27767716100682e+17, 1.27767716110682e+17, 1.277677161195884e+17, 1.27767716130682e+17, 1.27767716140682e+17, 1.27767716150682e+17, 1.277677161592758e+17, 1.27767716170682e+17, 1.27767716180682e+17, 1.277677161906821e+17, 1.277677161994319e+17, 1.27767716210682e+17, 1.27767716220682e+17, 1.27767716230682e+17, 1.277677162395882e+17, 1.27767716250682e+17, 1.27767716260682e+17, 1.27767716270682e+17, 1.277677162797445e+17, 1.27767716290682e+17, 1.27767716300682e+17, 1.27767716310682e+17, 1.277677163203695e+17, 1.27767716330682e+17, 1.27767716340682e+17, 1.27767716350682e+17, 1.277677163595882e+17, 1.27767716370682e+17, 1.27767716380682e+17, 1.27767716390682e+17, 1.277677164005257e+17, 1.27767716410682e+17, 1.27767716420682e+17, 1.27767716430682e+17, 1.277677164399008e+17, 1.277677164506821e+17, 1.27767716460682e+17, 1.27767716470682e+17, 1.277677164799008e+17, 1.27767716490682e+17, 1.27767716500682e+17, 1.27767716510682e+17, 1.277677165200571e+17, 1.27767716530682e+17, 1.27767716540682e+17, 1.27767716550682e+17, 1.277677165597445e+17, 1.27767716570682e+17, 1.27767716580682e+17, 1.27767716590682e+17, 1.27767716600057e+17, 1.27767716610682e+17, 1.27767716620682e+17, 1.27767716630682e+17, 1.277677166402132e+17, 1.27767716650682e+17, 1.27767716660682e+17, 1.27767716670682e+17, 1.277677166792758e+17, 1.27767716690682e+17, 1.27767716700682e+17, 1.277677167106821e+17, 1.277677167194319e+17, 1.27767716730682e+17, 1.27767716740682e+17, 1.27767716750682e+17, 1.277677167602132e+17, 1.27767716770682e+17, 1.27767716780682e+17, 1.27767716790682e+17, 1.277677167992758e+17, 1.27767716810682e+17, 1.27767716820682e+17, 1.27767716830682e+17, 1.277677168394321e+17, 1.27767716850682e+17, 1.27767716860682e+17, 1.27767716870682e+17, 1.277677168795884e+17, 1.27767716890682e+17, 1.27767716900682e+17, 1.27767716910682e+17, 1.277677169202132e+17, 1.27767716930682e+17, 1.27767716940682e+17, 1.27767716950682e+17, 1.277677169594319e+17, 1.27767716970682e+17, 1.27767716980682e+17, 1.27767716990682e+17, 1.277677169995882e+17, 1.27767717010682e+17, 1.27767717020682e+17, 1.27767717030682e+17, 1.277677170397444e+17, 1.27767717050682e+17, 1.27767717060682e+17, 1.27767717070682e+17, 1.277677170794321e+17, 1.27767717090682e+17, 1.27767717100682e+17, 1.27767717110682e+17, 1.277677171197445e+17, 1.27767717130682e+17, 1.27767717140682e+17, 1.27767717150682e+17, 1.277677171599008e+17, 1.27767717170682e+17, 1.27767717180682e+17, 1.27767717190682e+17, 1.27767717200057e+17, 1.27767717210682e+17, 1.27767717220682e+17, 1.27767717230682e+17, 1.27767717240057e+17, 1.27767717250682e+17, 1.27767717260682e+17, 1.27767717270682e+17, 1.277677172797445e+17, 1.27767717290682e+17, 1.27767717300682e+17, 1.27767717310682e+17, 1.277677173200571e+17, 1.27767717330682e+17, 1.277677173406821e+17, 1.27767717350682e+17, 1.277677173602132e+17, 1.27767717370682e+17, 1.27767717380682e+17, 1.27767717390682e+17, 1.277677173992758e+17, 1.27767717410682e+17, 1.27767717420682e+17, 1.27767717430682e+17, 1.27767717440057e+17, 1.27767717450682e+17, 1.27767717460682e+17, 1.27767717470682e+17, 1.277677174802131e+17, 1.27767717490682e+17, 1.27767717500682e+17, 1.27767717510682e+17, 1.277677175194321e+17, 1.27767717530682e+17, 1.27767717540682e+17, 1.27767717550682e+17, 1.277677175602132e+17, 1.27767717570682e+17, 1.27767717580682e+17, 1.27767717590682e+17, 1.277677176002132e+17, 1.27767717610682e+17, 1.27767717620682e+17, 1.27767717630682e+17, 1.277677176392756e+17, 1.27767717650682e+17, 1.27767717660682e+17, 1.27767717670682e+17, 1.277677176795882e+17, 1.27767717690682e+17, 1.27767717700682e+17, 1.27767717710682e+17, 1.277677177197445e+17, 1.27767717730682e+17, 1.27767717740682e+17, 1.27767717750682e+17, 1.277677177599008e+17, 1.27767717770682e+17, 1.27767717780682e+17, 1.27767717790682e+17, 1.277677177999008e+17, 1.27767717810682e+17, 1.27767717820682e+17, 1.27767717830682e+17, 1.277677178397445e+17, 1.27767717850682e+17, 1.27767717860682e+17, 1.27767717870682e+17, 1.277677178799008e+17, 1.27767717890682e+17, 1.27767717900682e+17, 1.27767717910682e+17, 1.27767717920057e+17, 1.27767717930682e+17, 1.27767717940682e+17, 1.27767717950682e+17, 1.27767717960682e+17, 1.27767717970682e+17, 1.27767717980682e+17, 1.27767717990682e+17, 1.27767718000682e+17, 1.27767718010682e+17, 1.27767718020682e+17, 1.27767718030682e+17, 1.277677180391195e+17, 1.277677180480257e+17, 1.27767718060682e+17, 1.27767718070682e+17, 1.27767718080682e+17, 1.27767718090682e+17, 1.27767718100682e+17, 1.277677181092758e+17, 1.277677181183383e+17, 1.27767718130682e+17, 1.27767718140682e+17, 1.277677181494321e+17, 1.27767718160682e+17, 1.27767718168182e+17, 1.27767718180682e+17, 1.277677181872445e+17, 1.27767718200682e+17, 1.27767718210682e+17, 1.277677182192758e+17, 1.277677182306821e+17, 1.277677182374008e+17, 1.277677182464634e+17, 1.27767718260682e+17, 1.27767718270682e+17, 1.277677182794319e+17, 1.27767718290682e+17, 1.277677182974007e+17, 1.277677183066195e+17, 1.27767718320682e+17, 1.27767718330682e+17, 1.277677183394321e+17},
			             {1.27767691700682e+17, 1.27767691710682e+17, 1.27767691720682e+17, 1.27767691730682e+17, 1.27767691740682e+17, 1.277676917506821e+17, 1.27767691760682e+17, 1.27767691770682e+17, 1.27767691780682e+17, 1.27767691790682e+17, 1.27767691800682e+17, 1.27767691810682e+17, 1.27767691820682e+17, 1.27767691830682e+17, 1.27767691840682e+17, 1.27767691850682e+17, 1.27767691860682e+17, 1.27767691870682e+17, 1.27767691880682e+17, 1.27767691890682e+17, 1.27767691900682e+17, 1.27767691910682e+17, 1.27767691920682e+17, 1.27767691930682e+17, 1.27767691940682e+17, 1.27767691950682e+17, 1.27767691960682e+17, 1.27767691970682e+17, 1.27767691980682e+17, 1.27767691990682e+17, 1.27767692000682e+17, 1.27767692010682e+17, 1.27767692020682e+17, 1.27767692030682e+17, 1.27767692040682e+17, 1.27767692050682e+17, 1.27767692060682e+17, 1.27767692070682e+17, 1.27767692080682e+17, 1.27767692090682e+17, 1.27767692100682e+17, 1.27767692110682e+17, 1.277676921206821e+17, 1.27767692130682e+17, 1.27767692140682e+17, 1.27767692150682e+17, 1.27767692160682e+17, 1.27767692170682e+17},
			             {1.27767692400682e+17, 1.27767692410682e+17, 1.27767692420682e+17, 1.27767692430682e+17, 1.27767692440682e+17, 1.27767692450682e+17, 1.27767692460682e+17, 1.27767692470682e+17, 1.27767692480682e+17, 1.27767692490682e+17, 1.27767692500682e+17, 1.27767692510682e+17, 1.27767692520682e+17, 1.27767692530682e+17, 1.27767692540682e+17, 1.27767692550682e+17, 1.27767692560682e+17, 1.27767692570682e+17, 1.27767692580682e+17, 1.27767692590682e+17, 1.27767692600682e+17, 1.27767692610682e+17},
			             {1.27767693370682e+17, 1.27767693380682e+17, 1.27767693390682e+17, 1.27767693400682e+17, 1.27767693410682e+17, 1.27767693420682e+17, 1.27767693430682e+17, 1.27767693440682e+17, 1.27767693450682e+17, 1.27767693460682e+17, 1.27767693470682e+17, 1.27767693480682e+17, 1.27767693490682e+17, 1.27767693500682e+17, 1.27767693510682e+17, 1.27767693520682e+17, 1.277676935306821e+17, 1.27767693540682e+17, 1.27767693550682e+17, 1.27767693560682e+17, 1.27767693570682e+17, 1.27767693580682e+17, 1.27767693590682e+17, 1.27767693600682e+17, 1.27767693610682e+17, 1.27767693620682e+17, 1.27767693630682e+17},
			             {1.27767691610682e+17, 1.27767691620682e+17, 1.27767691630682e+17, 1.27767691640682e+17, 1.27767691650682e+17, 1.27767691660682e+17, 1.27767691670682e+17, 1.27767691680682e+17, 1.27767691690682e+17, 1.27767691700682e+17, 1.27767691710682e+17, 1.27767691720682e+17, 1.27767691730682e+17, 1.27767691740682e+17, 1.277676917506821e+17, 1.27767691760682e+17, 1.27767691770682e+17, 1.27767691780682e+17, 1.27767691790682e+17, 1.27767691800682e+17, 1.27767691810682e+17, 1.27767691820682e+17, 1.27767691830682e+17, 1.27767691840682e+17, 1.27767691850682e+17, 1.27767691860682e+17, 1.27767691870682e+17, 1.27767691880682e+17, 1.27767691890682e+17, 1.27767691900682e+17, 1.27767691910682e+17, 1.27767691920682e+17, 1.27767691930682e+17, 1.27767691940682e+17, 1.27767691950682e+17, 1.27767691960682e+17, 1.27767691970682e+17, 1.27767691980682e+17, 1.27767691990682e+17, 1.27767692000682e+17, 1.27767692010682e+17, 1.27767692020682e+17, 1.27767692030682e+17, 1.27767692040682e+17, 1.27767692050682e+17, 1.27767692060682e+17, 1.27767692070682e+17, 1.27767692080682e+17, 1.27767692090682e+17, 1.27767692100682e+17, 1.27767692110682e+17, 1.277676921206821e+17, 1.27767692130682e+17, 1.27767692140682e+17, 1.27767692150682e+17, 1.27767692160682e+17, 1.27767692170682e+17, 1.27767692180682e+17, 1.27767692190682e+17, 1.27767692200682e+17, 1.27767692210682e+17, 1.27767692220682e+17, 1.27767692230682e+17, 1.27767692240682e+17, 1.27767692250682e+17, 1.27767692260682e+17, 1.27767692270682e+17, 1.27767692280682e+17, 1.27767692290682e+17, 1.27767692300682e+17, 1.27767692310682e+17, 1.27767692320682e+17, 1.27767692330682e+17, 1.27767692340682e+17, 1.27767692350682e+17, 1.27767692360682e+17, 1.27767692370682e+17},
			             {1.27767688240682e+17, 1.27767688250682e+17, 1.27767688260682e+17, 1.27767688270682e+17, 1.27767688280682e+17, 1.27767688290682e+17, 1.277676883006821e+17, 1.27767688310682e+17, 1.27767688320682e+17, 1.27767688330682e+17, 1.27767688340682e+17, 1.27767688350682e+17, 1.27767688360682e+17, 1.27767688370682e+17, 1.27767688380682e+17, 1.27767688390682e+17, 1.27767688400682e+17, 1.27767688410682e+17, 1.27767688420682e+17, 1.27767688430682e+17, 1.27767688440682e+17, 1.27767688450682e+17, 1.27767688460682e+17, 1.27767688470682e+17, 1.27767688480682e+17, 1.27767688490682e+17, 1.27767688500682e+17, 1.27767688510682e+17, 1.27767688520682e+17, 1.27767688530682e+17, 1.27767688540682e+17, 1.27767688550682e+17, 1.277676885606821e+17, 1.27767688570682e+17, 1.27767688580682e+17, 1.27767688590682e+17, 1.27767688600682e+17, 1.27767688610682e+17, 1.27767688620682e+17, 1.27767688630682e+17, 1.27767688640682e+17, 1.27767688650682e+17, 1.27767688660682e+17, 1.27767688670682e+17, 1.27767688680682e+17, 1.27767688690682e+17, 1.27767688700682e+17, 1.27767688710682e+17, 1.27767688720682e+17, 1.27767688730682e+17, 1.27767688740682e+17, 1.27767688750682e+17, 1.27767688760682e+17, 1.27767688770682e+17, 1.27767688780682e+17, 1.27767688790682e+17, 1.27767688800682e+17, 1.27767688810682e+17, 1.277676888206821e+17, 1.27767688830682e+17, 1.27767688840682e+17, 1.27767688850682e+17, 1.27767688860682e+17, 1.27767688870682e+17, 1.27767688880682e+17, 1.27767688890682e+17, 1.27767688900682e+17, 1.27767688910682e+17, 1.27767688920682e+17, 1.27767688930682e+17, 1.27767688940682e+17, 1.27767688950682e+17, 1.27767688960682e+17, 1.27767688970682e+17, 1.27767688980682e+17, 1.27767688990682e+17, 1.27767689000682e+17, 1.27767689010682e+17, 1.27767689020682e+17, 1.27767689030682e+17, 1.27767689040682e+17, 1.27767689050682e+17, 1.27767689060682e+17, 1.27767689070682e+17, 1.27767689080682e+17, 1.27767689090682e+17, 1.27767689100682e+17, 1.27767689110682e+17, 1.27767689120682e+17, 1.27767689130682e+17, 1.27767689140682e+17, 1.27767689150682e+17, 1.27767689160682e+17, 1.27767689170682e+17, 1.27767689180682e+17, 1.277676891906821e+17, 1.27767689200682e+17, 1.27767689210682e+17, 1.27767689220682e+17, 1.27767689230682e+17, 1.27767689240682e+17, 1.27767689250682e+17, 1.27767689260682e+17, 1.27767689270682e+17, 1.27767689280682e+17, 1.27767689290682e+17, 1.27767689300682e+17, 1.27767689310682e+17, 1.27767689320682e+17, 1.27767689330682e+17, 1.27767689340682e+17, 1.27767689350682e+17, 1.27767689360682e+17, 1.27767689370682e+17, 1.27767689380682e+17, 1.27767689390682e+17, 1.27767689400682e+17, 1.27767689410682e+17, 1.27767689420682e+17, 1.27767689430682e+17, 1.27767689440682e+17, 1.277676894506821e+17, 1.27767689460682e+17, 1.27767689470682e+17, 1.27767689480682e+17, 1.27767689490682e+17, 1.27767689500682e+17, 1.27767689510682e+17, 1.27767689520682e+17, 1.27767689530682e+17, 1.27767689540682e+17, 1.27767689550682e+17, 1.27767689560682e+17, 1.27767689570682e+17, 1.27767689580682e+17, 1.27767689590682e+17, 1.27767689600682e+17, 1.27767689610682e+17, 1.27767689620682e+17, 1.27767689630682e+17, 1.27767689640682e+17, 1.27767689650682e+17, 1.27767689660682e+17, 1.27767689670682e+17, 1.27767689680682e+17, 1.27767689690682e+17, 1.27767689700682e+17, 1.277676897106821e+17, 1.27767689720682e+17, 1.27767689730682e+17, 1.27767689740682e+17, 1.27767689750682e+17, 1.27767689760682e+17, 1.27767689770682e+17, 1.27767689780682e+17, 1.27767689790682e+17, 1.27767689800682e+17, 1.27767689810682e+17, 1.27767689820682e+17, 1.27767689830682e+17, 1.27767689840682e+17, 1.27767689850682e+17, 1.27767689860682e+17, 1.27767689870682e+17, 1.27767689880682e+17, 1.27767689890682e+17, 1.27767689900682e+17};
			mask_depths = {{187.6, 194.9}, {186.9, 195.7}, {185.0, 186.7, 195.9}, {184.9, 196.0}, {184.4, 196.1}, {181.5, 182.9, 196.6}, {177.2, 180.2, 196.9}, {176.4, 197.1}, {172.7, 197.1}, {172.4, 197.3}, {173.0, 197.6}, {176.5, 181.3, 197.8}, {183.0, 184.8, 190.9, 197.8}, {192.8, 196.8}}, {{184.7, 186.0}, {181.9, 183.2, 184.4, 186.5}, {181.9, 183.6, 184.6, 186.9}, {181.1, 183.9, 184.5, 187.0}, {181.1, 187.0}, {181.3, 187.2}, {181.3, 188.0}, {181.6, 189.0}, {181.9, 186.0, 189.2}, {186.9, 189.2}, {187.7, 188.7}}, {{179.6, 182.1}, {178.8, 182.5}, {178.8, 180.3, 185.6}, {181.0, 182.3, 185.6}, {184.4, 184.9}}, {{186.6, 190.6}, {186.7, 193.0, 195.8}, {187.2, 197.4}, {191.0, 198.1}, {198.2, 198.6}}, {{181.5, 185.2}, {180.1, 185.6}, {179.7, 179.8, 185.6, 185.7}, {179.5, 185.4}, {179.4, 185.3}, {179.3, 181.0, 185.0, 185.2}, {181.9, 184.6}}, {{168.7, 169.1}, {166.4, 169.6, 171.9}, {166.1, 172.4}, {166.1, 172.4}, {164.1, 164.5, 165.8, 172.1}, {163.4, 164.4, 165.3, 171.6}, {163.2, 164.7, 165.1, 171.8, 174.7}, {161.3, 177.6}, {159.4, 182.3}, {157.6, 182.6}, {157.2, 182.7}, {156.5, 182.8}, {155.5, 183.0}, {154.9, 183.0}, {153.0, 182.8}, {152.1, 182.1}, {150.8, 179.7, 181.0}, {150.4, 179.5}, {150.0, 179.3}, {149.7, 179.2}, {149.6, 179.6}, {149.4, 179.6}, {149.2, 179.7}, {148.8, 179.8}, {146.5, 181.9}, {146.2, 184.6}, {143.9, 185.2}, {143.5, 185.5}, {143.3, 185.5}, {142.9, 185.7}, {142.3, 185.7}, {141.9, 185.5}, {141.7, 185.3}, {141.5, 184.2}, {141.2, 183.8}, {141.0, 183.8}, {140.7, 183.7}, {140.3, 182.6}, {139.6, 182.4}, {139.0, 181.7}, {138.5, 181.5}, {137.9, 181.5}, {137.7, 181.7}, {136.7, 182.4}, {136.7, 183.4}, {136.8, 183.7}, {137.7, 183.8}, {138.1, 184.0}, {138.1, 184.2}, {138.2, 184.1}, {139.2, 184.1}, {139.3, 184.3}, {139.7, 184.2}, {140.3, 141.7, 184.3}, {141.8, 184.4}, {141.9, 184.7}, {142.0, 185.0}, {142.2, 185.4}, {142.3, 187.1}, {140.9, 187.4}, {141.0, 187.4}, {141.1, 187.5}, {141.0, 187.4}, {140.8, 187.1}, {140.1, 188.3}, {139.4, 188.7}, {138.8, 189.5}, {138.7, 189.8}, {138.6, 190.4}, {138.8, 191.0}, {137.8, 191.4}, {137.7, 191.4}, {137.2, 191.1}, {136.6, 190.9}, {134.5, 190.7}, {134.6, 189.1, 190.6}, {134.7, 189.0}, {134.8, 185.4, 188.1}, {134.7, 184.4}, {134.5, 184.2}, {134.4, 184.1}, {134.2, 184.1}, {134.0, 184.5}, {133.8, 184.9}, {133.5, 185.3}, {133.2, 185.7}, {132.9, 187.0}, {132.6, 186.9}, {132.3, 185.0, 186.8}, {131.9, 184.5}, {131.6, 183.9}, {131.4, 183.8}, {131.3, 183.7}, {131.2, 183.8}, {130.6, 184.9}, {130.7, 185.4}, {130.3, 177.9, 183.7, 185.0}, {130.7, 177.5, 184.2, 184.8}, {130.9, 177.1}, {130.9, 176.9}, {131.0, 177.8}, {131.4, 178.6}, {131.7, 179.1}, {131.9, 180.6}, {131.8, 180.7}, {131.8, 180.7}, {131.7, 181.1}, {131.8, 182.1}, {131.7, 182.2}, {131.5, 182.2}, {131.2, 182.1}, {131.1, 182.2}, {131.1, 182.5}, {131.4, 183.0}, {131.5, 183.3}, {131.2, 183.6}, {131.2, 183.6}, {131.1, 183.3}, {130.9, 183.1}, {130.8, 182.8}, {130.8, 181.1, 182.2}, {131.1, 181.0}, {131.4, 180.9}, {131.6, 181.0}, {131.8, 181.0}, {132.0, 180.8}, {131.7, 180.6}, {131.5, 180.4}, {131.5, 180.4}, {131.4, 180.0}, {131.6, 180.0}, {131.6, 179.9}, {131.6, 179.7}, {131.7, 179.8}, {131.9, 180.0}, {132.1, 179.7}, {132.4, 179.6}, {132.9, 179.3}, {132.5, 179.1}, {132.3, 179.3}, {132.6, 178.6, 179.6}, {133.0, 178.9}, {133.1, 178.8}, {133.7, 178.5}, {133.5, 177.9}, {133.3, 177.7}, {133.5, 177.9}, {133.9, 176.5, 178.1}, {134.2, 176.6}, {134.5, 173.8}, {134.9, 171.0}, {134.8, 170.5}, {134.8, 170.4}, {135.1, 170.4}, {135.2, 170.4}, {135.3, 168.7}, {135.4, 166.9, 168.2}, {135.6, 166.8}, {135.9, 166.9}, {136.7, 166.9}, {136.5, 166.5}, {136.5, 166.3}, {136.6, 166.4}, {136.8, 166.6}, {136.9, 166.9}, {136.8, 167.0}, {136.6, 169.1, 170.8}, {136.3, 172.2}, {136.4, 172.9}, {136.2, 173.1}, {136.2, 173.5}, {136.3, 173.6}, {136.4, 173.9}, {136.3, 173.6}, {136.3, 173.8}, {136.2, 173.8}, {135.9, 174.2}, {135.9, 174.3}, {135.6, 174.8}, {135.1, 174.8}, {135.1, 175.0}, {135.0, 175.0}, {134.8, 174.8}, {134.8, 174.4}, {134.7, 173.3}, {134.5, 173.1}, {134.5, 172.9}, {134.6, 172.6}, {134.5, 172.5}, {134.6, 169.8, 170.5, 172.4}, {135.2, 170.2, 171.3, 172.7}, {135.2, 170.2}, {135.5, 169.7}, {134.5, 169.7}, {133.8, 169.0}, {133.7, 168.3}, {134.2, 169.2}, {134.0, 169.0}, {134.2, 169.2}, {134.2, 169.2}, {134.2, 169.2}, {134.0, 169.0}, {134.0, 169.0}, {134.0, 169.0}, {134.1, 168.9}, {134.0, 168.6}, {133.9, 168.3}, {133.8, 168.2}, {134.0, 167.6}, {134.5, 168.0}, {134.7, 168.0}, {134.9, 168.0}, {135.0, 168.1}, {135.1, 168.2}, {135.1, 168.2}, {135.3, 168.2}, {135.9, 168.2}, {135.4, 167.6}, {135.4, 167.6}, {135.3, 166.4}, {136.2, 166.0, 167.1}, {136.0, 165.8}, {136.4, 166.7}, {136.4, 166.8}, {136.8, 166.8}, {136.9, 166.3}, {136.2, 166.1}, {136.1, 165.9}, {136.1, 165.5}, {136.2, 165.8}, {136.3, 166.2}, {136.0, 165.8}, {136.0, 165.8}, {136.1, 165.9}, {137.3, 167.0}, {136.7, 166.1}, {136.9, 166.3}, {136.2, 165.8}, {136.1, 165.7}, {136.1, 164.8}, {136.5, 165.8}, {136.5, 165.8}, {136.9, 166.2}, {136.8, 165.7}, {137.2, 165.9}, {137.1, 165.6}, {137.1, 165.6}, {137.4, 165.8}, {137.2, 165.7}, {137.4, 165.7}, {137.4, 165.7}, {137.7, 165.6}, {138.2, 165.7}, {138.3, 165.9}, {138.3, 166.1}, {138.3, 166.2}, {138.5, 166.4}, {138.3, 166.4}, {138.9, 167.2}, {138.9, 167.2}, {139.5, 167.4}, {138.9, 167.2}, {139.1, 167.4}, {138.8, 167.4}, {138.8, 167.4}, {138.7, 167.4}, {139.1, 167.8}, {138.8, 167.8}, {139.0, 168.2}, {138.8, 168.4}, {138.4, 168.4}, {138.4, 168.6}, {137.9, 168.7}, {137.9, 169.2}, {137.8, 169.1}, {138.1, 169.5}, {137.9, 169.5}, {138.1, 169.9}, {138.1, 169.9}, {138.0, 169.9}, {137.6, 169.9}, {137.6, 170.1}, {137.6, 170.3}, {137.6, 170.3}, {137.6, 170.1}, {137.6, 170.1}, {137.4, 169.9}, {137.3, 170.0}, {137.4, 170.3}, {137.2, 170.3}, {137.3, 170.6}, {137.3, 170.8}, {137.6, 170.9, 172.0}, {137.1, 172.1, 174.2, 174.8}, {137.3, 172.3, 174.0, 175.0}, {137.1, 172.2, 173.8, 174.7}, {137.1, 172.2, 173.8, 174.7}, {137.2, 172.8, 173.9, 174.5}, {137.7, 175.4}, {137.7, 175.4}, {137.7, 175.4}, {138.0, 175.5}, {137.8, 175.5}, {138.0, 175.7}, {140.1, 175.9}, {140.5, 176.1}, {140.9, 176.3}, {141.4, 176.2}, {143.5, 176.3}, {144.2, 176.5}, {144.2, 176.5}, {144.2, 176.5}, {144.6, 176.9}, {144.4, 176.9}, {145.0, 177.7, 180.7}, {146.1, 181.4}, {145.1, 181.4}, {145.5, 181.6}, {144.8, 181.3}, {144.8, 181.3}, {144.8, 180.7}, {145.0, 181.1}, {144.8, 180.9}, {145.0, 181.1}, {145.4, 182.1}, {145.4, 182.3}, {146.5, 182.4}, {147.0, 182.6}, {145.7, 182.4}, {145.7, 182.4}, {145.7, 181.3}, {146.0, 182.7}, {146.0, 182.7}, {146.2, 182.9}, {145.9, 182.6}, {146.1, 147.1, 182.8}, {147.2, 183.0}, {147.4, 183.1}, {147.6, 183.4}, {147.5, 183.2}, {147.7, 183.6}, {147.4, 183.4}, {147.3, 183.3}, {148.0, 183.5}, {147.8, 183.3}, {148.2, 183.7}, {148.2, 183.8}, {148.4, 183.8}, {148.1, 183.3}, {148.3, 183.5}, {148.4, 183.4}, {147.8, 183.1}, {147.8, 183.1}, {148.4, 183.4}, {148.2, 182.8}, {148.5, 183.3}, {149.2, 184.0}, {149.7, 184.0}, {148.9, 183.1}, {149.1, 183.5}, {148.7, 183.1}, {148.6, 183.2}, {149.2, 184.0}, {149.2, 184.0}, {149.3, 184.1}, {149.3, 183.9}, {149.5, 183.9}, {149.5, 184.0}, {149.5, 183.8}, {149.7, 184.1}, {150.0, 184.4}, {150.2, 184.4}, {149.8, 184.1}, {150.0, 184.2}, {149.6, 184.0}, {149.4, 183.8}, {149.9, 184.3}, {149.7, 183.4}, {150.0, 183.7}, {150.2, 183.9}, {151.2, 184.1}, {150.0, 183.7}, {150.0, 184.0}, {149.9, 183.9}, {150.5, 184.7}, {150.5, 184.5}, {150.9, 184.9}, {152.1, 184.8}, {151.4, 183.2}, {151.8, 183.0}, {151.5, 182.5}, {151.5, 182.5}, {151.9, 182.7}, {151.8, 182.5}, {151.8, 182.8}, {151.8, 182.8}, {151.7, 182.8}, {151.7, 182.8}, {151.9, 183.0}, {151.8, 182.9}, {151.8, 182.9}, {152.0, 183.2}, {152.4, 183.4}, {151.7, 182.9}, {151.7, 183.1}, {151.0, 182.5}, {151.6, 183.3}, {151.4, 182.5}, {151.0, 183.9, 187.3, 188.7}, {151.0, 183.9, 187.1, 188.9}, {152.0, 184.1, 187.0, 189.3}, {150.8, 183.5, 185.0, 189.0}, {151.0, 183.6, 184.8, 189.4}, {150.4, 183.2, 184.0, 189.2}, {150.4, 189.4}, {150.5, 189.5}, {150.7, 189.9}, {150.5, 189.7}, {150.4, 189.8}, {150.5, 190.0}, {150.1, 189.8}, {150.2, 190.1}, {150.2, 190.1}, {150.2, 190.1}, {150.8, 182.9, 185.4, 190.0}, {149.6, 181.4, 185.8, 187.1}, {149.6, 181.4}, {149.6, 181.4}, {149.7, 181.6}, {149.5, 181.4}, {149.7, 181.7}, {149.7, 181.5}, {150.2, 181.2}, {149.7, 180.1}, {149.9, 180.1}, {149.3, 179.3}, {149.3, 179.3}, {149.3, 179.3}, {149.3, 179.5}, {149.3, 179.5}, {149.3, 179.3}, {149.1, 178.6}, {149.0, 177.1}, {148.8, 176.1}, {149.2, 176.8}, {149.2, 176.8}, {149.2, 176.9}, {148.3, 176.4}, {148.3, 176.4}, {148.3, 176.4}, {148.3, 176.5}, {148.1, 176.4}, {147.9, 175.8}, {147.8, 175.9}, {147.6, 175.7}, {147.5, 175.8}, {147.4, 175.9}, {147.4, 175.9}, {147.4, 175.7}, {147.6, 175.9}, {147.2, 175.7}, {146.7, 175.2}, {146.7, 175.0}, {146.9, 175.6}, {146.7, 175.4}, {147.1, 175.6}, {147.1, 175.5}, {147.2, 175.5}, {147.8, 175.6}, {147.5, 175.2}, {147.9, 175.2}, {147.9, 174.9}, {148.0, 174.0}, {148.9, 174.5}, {148.7, 174.3}, {149.3, 174.9}, {149.3, 174.9}, {149.8, 175.0}, {149.2, 175.6}, {149.6, 175.8}, {149.1, 175.3}, {149.1, 175.3}, {149.3, 175.1}, {149.6, 175.4}, {149.2, 175.4}, {149.2, 175.4}, {148.9, 175.3}, {149.2, 175.8}, {149.2, 175.8}, {148.8, 175.3}, {149.3, 175.3}, {148.7, 174.5}, {148.1, 173.9}, {147.9, 173.1}, {147.9, 172.0, 172.6, 174.5}, {147.5, 170.9, 172.8, 173.5}, {148.5, 172.0}, {148.5, 172.0}, {147.5, 171.2}, {148.3, 171.4}, {147.5, 171.2}, {146.9, 171.0}, {147.2, 171.3}, {147.2, 170.9}, {147.1, 170.4}, {147.2, 171.8}, {147.2, 170.9}, {146.9, 170.6}, {147.6, 170.6}, {147.7, 169.5}, {146.7, 169.1}, {146.3, 168.7}, {146.3, 167.3, 168.3}, {146.6, 166.9}, {146.6, 167.8}, {146.4, 167.6}, {146.6, 167.9}, {146.6, 167.9}, {147.1, 167.8}, {146.4, 166.6}, {147.0, 166.6}, {146.0, 165.7}, {146.0, 165.7}, {145.9, 164.5}, {146.2, 165.7}, {145.8, 165.5}, {146.3, 166.2}, {146.4, 166.5}, {145.9, 165.7}, {146.4, 166.3}, {145.6, 166.1}, {145.6, 166.1}, {145.6, 166.1}, {145.3, 165.4}, {145.7, 165.8}, {145.3, 165.6}, {145.9, 166.3}, {145.9, 166.3}, {145.6, 166.3}, {146.4, 166.4}, {145.4, 166.6, 167.6}, {145.4, 167.8}, {145.0, 167.4}, {145.1, 166.5}, {145.7, 166.7}, {145.3, 166.7}, {145.8, 167.2}, {145.8, 167.2}, {145.1, 166.7}, {145.1, 166.9}, {144.9, 166.8}, {144.7, 166.9}, {144.7, 167.1}, {144.5, 167.1}, {144.4, 167.0}, {144.3, 167.1}, {144.1, 166.9}, {144.2, 166.9}, {144.2, 167.1}, {144.2, 167.1}, {144.1, 167.1}, {144.1, 166.9}, {144.1, 166.9}, {144.4, 167.0}, {144.5, 166.9}, {144.7, 166.9}, {144.6, 167.0}, {144.6, 167.0}, {144.7, 167.1}, {144.7, 167.1}, {144.9, 167.3}, {144.9, 167.3}, {145.1, 167.5}, {145.5, 167.8}, {146.1, 168.1}, {145.5, 168.6, 169.6, 170.2}, {145.7, 168.8, 169.4, 170.4}, {145.4, 170.2}, {145.1, 170.0}, {146.0, 171.0}, {145.6, 171.0}, {146.1, 171.9}, {146.3, 172.5}, {146.9, 172.7}, {147.3, 172.9}, {146.0, 172.0}, {146.0, 172.0}, {146.9, 172.7}, {146.5, 172.7}, {147.2, 173.8}, {147.2, 174.2}, {147.4, 174.4}, {147.6, 174.8}, {147.4, 174.5}, {147.6, 174.5}, {147.5, 174.4}, {147.7, 174.6}, {147.7, 174.6}, {148.2, 175.3}, {149.3, 176.4}, {148.5, 176.6}, {149.1, 176.6}, {149.1, 176.6}, {149.0, 176.3}, {149.0, 176.1}, {149.2, 176.7}, {149.8, 177.4}, {149.5, 177.4}, {150.3, 178.7, 181.4, 182.2}, {151.4, 178.9, 180.1, 182.4, 183.3, 183.7}, {151.5, 179.0, 179.6, 182.4, 183.0, 183.8}, {151.5, 183.8}, {151.9, 184.4}, {152.3, 184.8}, {152.6, 185.1}, {153.2, 186.1}, {153.6, 186.3}, {153.7, 186.2}, {153.4, 185.9}, {153.4, 185.9}, {153.3, 186.0}, {154.0, 187.0}, {154.0, 187.2}, {154.4, 189.0}, {155.2, 189.2}, {155.3, 188.9}, {155.5, 188.9}, {155.5, 188.4}, {156.4, 189.1}, {156.6, 189.1}, {157.0, 189.1}, {157.0, 188.9}, {157.2, 189.0}, {157.4, 189.0}, {158.2, 189.1}, {157.9, 188.9}, {158.1, 189.1}, {158.0, 189.0}, {158.3, 189.4}, {158.8, 190.2}, {158.8, 190.2}, {159.4, 190.4}, {158.8, 189.8}, {158.8, 190.0}, {158.8, 190.0}, {158.5, 189.6}, {158.6, 189.8}, {158.4, 189.6}, {158.3, 189.9}, {158.3, 190.1}, {158.0, 189.7}, {157.8, 189.3}, {157.4, 187.4, 188.2, 189.5}, {157.0, 187.2, 188.6, 189.2}, {157.0, 187.6}, {156.9, 187.5}, {157.2, 187.1}, {156.3, 187.0}, {156.3, 187.0}, {156.0, 186.8}, {156.2, 187.4}, {156.0, 187.0}, {155.9, 187.4}, {156.2, 187.5}, {156.4, 187.6}, {155.7, 186.6}, {155.7, 186.6}, {155.2, 186.0}, {155.2, 185.8}, {155.6, 186.2}, {155.6, 186.2}, {155.7, 186.1}, {155.4, 185.4}, {154.9, 184.8}, {154.9, 184.6}, {154.8, 184.5}, {154.3, 185.4}, {154.1, 185.4}, {154.0, 185.4}, {154.6, 185.6}, {153.5, 184.9}, {153.5, 184.9}, {153.1, 184.2}, {153.1, 183.9}, {153.2, 183.6}, {153.3, 184.1}, {153.2, 183.9}, {153.0, 183.8}, {153.0, 183.8}, {153.3, 183.8}, {153.4, 183.8}, {153.2, 183.6}, {153.4, 183.8}, {153.3, 183.7}, {153.2, 183.6}, {153.3, 183.5}, {153.7, 183.7}, {154.3, 183.5}, {154.9, 183.8}, {155.1, 183.6}, {155.4, 156.5, 183.5}, {157.1, 183.3}, {157.2, 183.0}, {157.6, 183.0}, {157.8, 182.8}, {158.2, 182.8}, {158.3, 183.0}, {158.4, 183.0}, {158.4, 183.2}, {158.4, 183.5}, {158.5, 183.7}, {158.5, 183.7}, {158.5, 183.7}, {158.3, 183.7}, {158.6, 183.9}, {158.6, 184.1}, {158.8, 184.2}, {158.7, 184.3}, {158.6, 184.6}, {158.9, 185.1}, {158.9, 185.1}, {159.3, 185.3}, {159.2, 185.2}, {159.2, 185.2}, {159.2, 185.2}, {159.4, 185.4}, {159.8, 185.6}, {160.2, 185.6}, {160.3, 185.5}, {160.5, 185.7}, {160.4, 185.7}, {160.4, 185.6}, {160.7, 186.0}, {160.5, 185.8}, {160.8, 186.1}, {161.1, 186.2}, {161.2, 186.0}, {161.0, 185.9}, {160.5, 185.4}, {160.5, 185.4}, {160.6, 185.5}, {160.9, 185.7}, {160.8, 186.2}, {160.8, 185.6}, {160.8, 185.6}, {160.6, 185.5}, {160.6, 185.3}, {160.4, 185.1}, {160.4, 185.4}, {159.9, 185.5}, {159.6, 185.7}, {160.2, 186.6}, {159.8, 186.6}, {159.3, 185.4, 186.0, 187.0}, {159.2, 185.6, 186.5, 187.1}, {159.2, 185.6}, {159.1, 185.3}, {158.5, 184.5}, {158.5, 184.3}, {158.3, 183.9}, {158.3, 183.8}, {158.1, 183.8}, {158.1, 183.8}, {158.1, 183.9}, {157.9, 183.9}, {157.9, 182.7, 183.3, 184.1}, {157.7, 182.5, 183.5, 183.9}, {157.4, 182.7}, {157.4, 182.8}, {157.3, 182.7}, {157.1, 182.3}, {156.9, 182.2}, {156.5, 181.7}, {156.5, 181.7}, {156.0, 181.3}, {156.3, 181.5}, {156.1, 181.2}, {156.0, 180.9}, {156.0, 181.0}, {156.0, 179.9}, {156.0, 179.9}, {156.4, 179.5}, {156.3, 178.7}, {155.6, 178.5}, {154.7, 177.9}, {154.7, 177.9}, {155.1, 176.7}, {155.2, 178.2}, {154.8, 178.0}, {155.3, 178.8}, {155.5, 179.0}, {156.5, 178.7}, {154.8, 178.9}, {154.8, 178.9}, {154.1, 178.0}, {154.8, 178.3}, {154.6, 177.6}, {154.9, 178.2}, {154.7, 178.7}, {154.4, 178.9}, {154.1, 180.9}, {153.9, 180.8}, {153.9, 180.8}, {154.1, 181.0}, {154.2, 181.0}, {154.4, 181.0}, {154.0, 182.5}, {154.0, 183.3}, {153.9, 183.1}, {154.0, 183.0}, {154.1, 182.0}, {154.0, 182.9}, {153.8, 182.9}, {154.0, 183.1}, {154.0, 183.0}, {154.4, 183.1}, {153.7, 183.2}, {153.7, 183.4}, {153.6, 183.2}, {153.5, 183.2}, {153.3, 183.0}, {153.4, 182.6}, {153.3, 183.7}, {153.3, 183.7}, {154.6, 184.2}, {154.3, 157.4, 184.0}, {159.5, 184.4}, {158.3, 184.1}, {158.3, 184.1}, {158.3, 183.8}, {158.3, 183.8}, {158.1, 184.1}, {158.4, 184.4}, {158.4, 184.4}, {158.6, 184.6}, {158.4, 184.8}, {158.6, 184.9}, {158.6, 185.9}, {158.4, 185.9}, {158.0, 185.8}, {157.8, 185.5}, {157.8, 185.7}, {157.6, 185.6}, {158.0, 186.4}, {158.0, 186.4}, {158.2, 186.5}, {158.6, 187.9}, {158.6, 187.7}, {158.2, 187.2}, {158.2, 187.0, 187.8, 188.2}, {158.0, 186.9, 187.6, 188.0}, {158.2, 187.0, 187.8, 188.2}, {158.2, 187.0, 187.8, 188.0}, {158.5, 188.2}, {158.7, 188.1}, {158.7, 188.1}, {158.6, 188.0}, {159.1, 188.3}, {159.1, 188.2}, {159.5, 188.3}, {159.5, 188.1}, {160.0, 188.0}, {160.0, 187.4}, {159.4, 186.9}, {159.0, 186.5}, {159.6, 187.0}, {159.4, 186.8}, {159.8, 187.3}, {160.2, 187.8}, {161.1, 187.8}, {161.2, 188.0}, {161.2, 187.9}, {161.3, 188.1}, {161.6, 188.0}, {160.9, 187.5}, {160.9, 187.5}, {160.8, 186.3}, {161.0, 186.3}, {161.4, 186.6}, {161.4, 186.6}, {161.4, 186.9}, {161.6, 187.2}, {161.7, 187.7}, {162.5, 188.3}, {162.7, 188.3}, {163.7, 187.8}, {163.4, 187.9}, {162.1, 187.4}, {161.6, 186.8}, {162.0, 184.3}, {162.0, 186.9}, {161.7, 186.7}, {162.5, 187.3}, {162.3, 187.2}, {164.6, 187.4}, {163.8, 187.9}, {164.6, 188.3}, {164.0, 188.1}, {163.5, 187.6}, {163.1, 185.5}, {163.6, 186.9}, {163.4, 186.5}, {163.2, 186.3}, {161.9, 187.1}, {162.2, 188.0}, {161.7, 188.9}, {162.7, 190.0}, {162.8, 190.3}, {162.5, 190.4}, {162.2, 189.9}, {162.4, 190.1}, {162.4, 189.0}, {163.2, 189.2}, {163.4, 190.2}, {163.7, 191.2}, {163.6, 191.1}, {164.2, 191.3}, {164.4, 191.4}, {163.6, 191.1}, {163.2, 190.9}, {163.4, 191.1}, {163.2, 191.3}, {163.3, 191.8}, {163.4, 192.4}, {163.6, 193.4}, {163.4, 193.4}, {163.7, 193.7}, {163.7, 193.9}, {163.4, 193.7}, {163.8, 193.8}, {163.4, 194.0}, {163.0, 194.7}, {163.0, 194.7}, {163.4, 195.1}, {163.2, 195.0}, {163.7, 195.4}, {163.9, 195.7}, {165.1, 195.7}, {165.0, 195.2}, {165.2, 195.2}, {166.3, 195.3}, {167.0, 195.3}, {168.2, 169.4, 195.6}, {169.5, 195.7}, {170.8, 196.0}, {170.9, 196.1}, {171.9, 196.1}, {172.2, 196.3}, {172.5, 196.6}, {172.9, 196.6}, {172.8, 196.5}, {173.8, 196.7}, {174.0, 196.7}, {173.9, 196.5}, {174.1, 196.5}, {174.2, 196.6}, {174.2, 196.6}, {174.1, 196.5}, {173.6, 196.4}, {173.1, 196.6}, {172.6, 196.3}, {172.6, 196.5}, {172.4, 196.0}, {172.5, 195.8}, {172.8, 196.9}, {172.8, 196.9}, {173.3, 198.7}, {173.2, 198.9}, {172.4, 198.7}, {171.9, 198.3}, {172.5, 198.7}, {172.3, 198.1}, {172.6, 199.2}, {172.6, 199.2}, {172.9, 199.5, 201.0}, {173.6, 201.1}, {173.5, 201.4, 203.0}, {173.7, 203.3}, {173.8, 203.2}, {173.7, 203.7}, {173.4, 203.4}, {173.4, 203.0}, {173.9, 203.5}, {173.7, 203.3}, {174.0, 203.7}, {174.2, 203.8}, {174.2, 203.8}, {174.1, 203.7}, {173.5, 203.3, 204.2, 204.8}, {173.5, 203.5, 204.2, 204.8}, {173.5, 203.7, 204.1, 204.9}, {174.1, 205.3}, {174.3, 205.1}, {174.6, 205.0}, {174.7, 204.3}, {174.6, 203.8}, {174.2, 203.4}, {174.2, 203.3}, {174.2, 202.5}, {174.6, 202.5}, {174.4, 202.3}, {174.7, 202.4}, {175.1, 202.7}, {175.1, 202.7, 203.8}, {174.9, 203.9}, {174.6, 203.9}, {174.6, 203.9}, {174.7, 204.0}, {174.8, 203.9}, {174.6, 203.6}, {174.4, 203.2}, {174.9, 203.6}, {174.5, 203.4}, {175.1, 204.1}, {175.1, 204.3}, {174.9, 204.4}, {174.7, 204.7}, {174.7, 204.7}, {175.1, 204.9}, {174.4, 205.0}, {174.4, 205.0}, {174.1, 204.5}, {174.8, 203.9, 204.8}, {174.8, 203.7}, {175.6, 204.5}, {176.2, 205.0}, {176.6, 205.3}, {177.6, 205.3}, {176.8, 205.5}, {177.6, 205.7}, {177.1, 205.0}, {176.8, 203.6}, {176.8, 202.6}, {177.5, 202.7}, {177.3, 202.7}, {177.6, 203.0}, {177.9, 203.3}, {178.1, 203.6}, {178.1, 203.7}, {178.2, 203.8}, {178.5, 203.9}, {179.7, 204.0}, {179.3, 203.5}, {179.5, 203.5}, {179.1, 202.8}, {180.0, 202.5}, {179.8, 202.3}, {180.6, 202.9}, {180.6, 202.9}, {180.7, 202.9}, {181.3, 203.0}, {181.2, 203.0}, {181.6, 204.1}, {181.6, 204.3}, {181.6, 204.4}, {182.2, 204.6}, {181.8, 205.0}, {181.4, 204.5}, {181.1, 203.3}, {181.8, 204.1}, {181.4, 204.0}, {181.4, 204.2}, {181.3, 204.4}, {181.2, 204.4}, {180.7, 204.2}, {181.0, 204.4}, {180.5, 203.7}, {180.1, 203.2, 204.8}, {180.4, 205.1}, {180.3, 204.7}, {180.5, 204.6}, {180.1, 205.4}, {180.1, 205.2}, {180.3, 204.9}, {179.4, 203.6}, {179.4, 203.6}, {179.2, 203.3}, {179.2, 203.1}, {179.1, 203.0}, {178.9, 203.0}, {178.8, 202.9}, {178.7, 202.8}, {178.5, 202.8}, {178.7, 203.1}, {178.7, 203.1}, {178.5, 203.2}, {178.1, 201.4, 202.6}, {178.1, 201.2}, {178.0, 201.0}, {178.0, 200.7}, {177.9, 200.8}, {177.8, 201.3}, {177.8, 201.3}, {177.7, 201.4}, {177.7, 201.4}, {177.5, 201.4}, {177.4, 201.3}, {177.4, 201.3}, {177.2, 201.1}, {177.0, 200.7}, {177.1, 200.8}, {176.9, 200.6}, {177.1, 200.8}, {176.9, 201.0}, {177.0, 201.1}, {177.0, 201.1}, {176.8, 200.9}, {176.5, 201.2}, {176.0, 201.3}, {176.0, 201.8}, {176.1, 201.9}, {176.4, 202.4}, {176.1, 202.1}, {176.2, 202.0}, {176.3, 200.4, 201.2, 202.2}, {176.1, 200.2, 201.3, 201.7}, {176.3, 200.2}, {176.5, 199.8}, {176.0, 200.1}, {175.6, 199.9}, {175.6, 199.9}, {175.7, 199.6}, {175.9, 200.1}, {176.2, 200.5}, {176.2, 200.5}, {176.4, 199.9}, {176.2, 199.3}, {176.1, 198.8}, {176.0, 198.2}}, {{134.2, 140.2}, {132.2, 133.5, 140.9, 141.2}, {131.9, 141.2, 142.5}, {131.0, 131.6, 143.3}, {128.7, 130.0, 144.1, 144.4}, {127.1, 144.6}, {125.9, 143.6}, {124.3, 124.9, 141.2, 142.1}, {121.7, 123.0, 141.0}, {121.5, 141.1}, {121.1, 121.4, 141.3, 141.5}, {121.1, 141.6}, {121.1, 141.4}, {121.1, 140.9}, {121.1, 140.9}, {121.1, 141.4}, {120.9, 142.7}, {120.7, 143.3}, {120.4, 144.5}, {120.4, 145.4}, {120.1, 120.4, 146.3, 147.3}, {120.1, 147.1, 147.2}, {120.1, 121.4, 148.4}, {121.7, 148.8}, {122.0, 122.3, 148.4, 149.2}, {122.3, 122.7, 149.6}, {123.1, 149.9}, {123.6, 150.2}, {124.6, 149.9}, {125.9, 149.8}, {125.9, 149.6, 151.1, 151.5}, {126.8, 150.1, 150.8, 151.6}, {127.1, 151.7}, {127.4, 127.8, 151.8, 151.9}, {127.8, 152.2}, {128.1, 128.4, 146.9, 147.7, 150.8, 151.5, 152.5}, {128.7, 129.7, 146.9, 148.1, 150.8, 151.7, 152.7}, {130.3, 130.6, 146.7, 147.9, 150.6, 151.7, 152.7}, {130.6, 146.5, 147.2, 149.9, 151.6, 152.2}, {131.0, 131.3, 146.3, 146.8, 149.3}, {130.3, 146.3, 147.5, 149.0}, {131.0, 131.6, 146.0, 148.1, 148.7}, {132.2, 133.5, 146.6, 146.8}, {133.7, 133.8, 146.9, 147.1}, {134.3, 147.1}, {134.8, 136.1, 146.4, 147.1}, {136.4, 146.4}, {136.7, 146.3}}, {{120.7, 124.9}, {119.0, 126.7, 128.0}, {118.5, 129.9}, {117.9, 130.7}, {117.5, 130.7}, {116.1, 132.0}, {114.8, 133.4}, {114.2, 135.2, 136.4}, {113.6, 138.5}, {112.7, 139.7}, {112.5, 140.6}, {112.4, 141.6}, {112.8, 142.2}, {114.0, 142.5}, {115.3, 143.8}, {114.8, 143.5}, {115.0, 143.9}, {115.7, 144.6}, {116.5, 142.1}, {116.8, 141.6}, {118.7, 140.7}, {130.9, 133.4}}, {{125.0, 126.0}, {118.1, 118.6, 124.8, 127.4, 130.7, 131.3}, {112.6, 115.7, 120.8, 121.6, 128.7, 129.2, 131.9, 134.8}, {107.9, 135.5}, {107.4, 129.6, 130.5, 135.7}, {107.3, 129.5, 133.9, 135.8}, {107.3, 129.7}, {107.4, 130.0, 147.6, 149.5}, {107.3, 130.1, 147.5, 150.5}, {107.0, 129.8, 146.6, 150.4}, {107.3, 130.6, 146.1, 150.3}, {107.8, 131.1, 145.6, 151.0, 153.7}, {109.2, 131.8, 145.1, 153.6}, {109.8, 134.2, 143.4, 153.9, 155.6}, {111.2, 157.9}, {112.5, 160.7}, {114.3, 115.8, 161.5}, {117.0, 164.8}, {119.5, 164.8}, {120.9, 164.5}, {122.2, 164.1}, {123.2, 159.9, 161.3, 164.0}, {123.7, 158.1, 159.7, 161.8, 164.2}, {125.6, 126.9, 157.1, 162.1, 164.6, 165.7}, {130.5, 152.5, 162.1, 165.9}, {133.8, 150.6, 162.1, 166.3}, {135.7, 139.3, 162.4, 165.9}}, {{137.3, 137.9}, {136.9, 138.7}, {126.6, 128.9, 140.6, 142.9}, {124.6, 143.4}, {120.6, 123.6, 143.7, 149.6, 150.2}, {119.9, 146.1, 149.6, 150.5}, {114.8, 115.3, 117.6, 118.2, 119.7, 151.3}, {114.4, 115.7, 117.0, 118.6, 119.2, 135.8, 142.8, 153.0}, {114.0, 127.8, 135.1, 142.8, 152.8}, {113.7, 126.5, 127.4, 142.8, 143.1, 152.5}, {112.5, 125.9, 126.2, 143.1, 144.4, 151.5}, {112.3, 124.9, 125.5, 144.7, 145.0, 151.1}, {111.4, 124.3, 124.6, 145.0, 149.1}, {110.7, 123.9, 124.3, 145.0, 148.0}, {110.6, 123.0, 123.9}, {109.8, 121.7, 122.7}, {108.6, 121.4, 121.7}, {107.6, 121.1, 121.4}, {106.7, 120.4, 121.1}, {106.2, 119.1, 120.4}, {105.1, 118.5, 118.8}, {105.1, 117.9, 118.2}, {105.0, 117.9}, {104.7, 117.2, 117.5}, {104.1, 117.2}, {103.8, 117.2}, {103.6, 117.2}, {103.6, 117.2}, {103.5, 117.2}, {103.5, 117.2}, {103.8, 117.2}, {103.2, 117.5}, {102.7, 117.9, 118.2}, {103.0, 118.2, 119.5}, {102.6, 119.5}, {105.1, 119.5, 120.1}, {107.0, 120.4, 121.1}, {109.8, 121.4, 122.0}, {111.3, 122.3, 123.0}, {111.8, 123.0, 123.3}, {111.8, 123.6}, {111.5, 123.6, 123.9}, {111.6, 124.3, 124.9}, {111.7, 125.2, 125.5}, {111.7, 125.5, 125.9}, {109.5, 125.9, 126.2}, {109.2, 126.5, 127.1}, {109.0, 127.1}, {108.8, 127.1}, {109.1, 127.1, 127.8}, {108.9, 127.8}, {109.0, 128.1, 129.4}, {109.5, 130.0, 130.6}, {110.0, 130.6, 131.0}, {110.4, 131.3, 132.4}, {111.1, 132.9}, {110.8, 132.9, 133.2}, {109.9, 133.5, 134.8}, {110.0, 135.1, 135.8}, {110.8, 136.1, 146.8}, {110.5, 148.2}, {110.6, 149.0}, {110.4, 149.0}, {110.6, 148.7}, {110.5, 148.3}, {111.4, 147.6}, {111.4, 147.6}, {111.9, 147.8}, {112.4, 148.0}, {111.2, 148.1}, {111.6, 145.6, 146.2, 148.3}, {112.3, 145.3, 146.7, 148.0}, {116.3, 145.5, 147.1, 148.4}, {117.3, 120.1, 145.6, 147.3, 148.6}, {123.3, 143.6, 146.8, 148.2}, {124.6, 128.1, 129.2, 135.7, 140.5, 142.2, 146.8, 147.2}, {127.7, 128.1, 135.7, 136.8}}, {{103.7, 104.7}, {103.9, 105.7, 108.1, 108.5}, {104.1, 107.8, 108.4, 108.7}, {104.8, 107.5, 110.5, 112.6}, {104.4, 106.4, 109.2, 112.7, 116.9, 118.8}, {104.2, 105.7, 107.2, 112.2, 116.0, 118.1}, {105.5, 106.2, 107.0, 112.5, 116.2, 117.7}, {106.6, 112.2, 117.1, 118.5}, {107.8, 113.0, 117.8, 119.3}, {108.3, 113.3, 117.9, 119.6}, {108.2, 113.4, 117.8, 119.7}, {107.9, 113.6, 117.3, 119.7, 131.4, 132.2}, {107.5, 115.0, 116.7, 119.4, 130.3, 131.8}, {107.3, 108.1, 109.4, 118.8, 123.6, 124.0, 129.9, 131.0}, {107.1, 107.5, 109.6, 117.1, 122.8, 123.6, 129.5, 130.7}, {109.6, 116.7, 122.1, 123.2, 129.3, 130.5}, {109.8, 116.7, 121.7, 122.6, 129.1, 130.5}, {110.6, 117.3, 121.9, 123.2, 129.0, 131.3}, {111.6, 118.2, 121.1, 124.2, 128.4, 129.3, 133.2}, {109.2, 111.1, 112.1, 129.1, 129.7, 133.9}, {108.8, 110.9, 111.7, 134.3}, {107.7, 134.7}, {107.0, 134.2}, {106.6, 134.5}, {103.8, 104.4, 105.9, 134.9}, {101.6, 103.5, 104.8, 105.6, 135.4, 136.4}, {101.2, 136.5}, {100.5, 134.3, 136.4}, {99.7, 132.4, 133.9}, {99.7, 132.4}, {99.8, 131.2}, {99.7, 130.7}, {102.7, 130.6}, {103.0, 104.9, 130.6}, {104.8, 130.8}, {104.4, 131.1, 133.6}, {104.0, 133.8}, {102.5, 134.5}, {101.7, 134.8}, {101.7, 134.5}, {101.7, 134.5}, {101.6, 134.5}, {101.2, 133.9}, {101.0, 132.4}, {100.9, 132.5}, {99.1, 100.6, 132.2}, {99.1, 132.2}, {99.3, 132.8}, {99.4, 132.5}, {99.3, 132.4}, {99.6, 132.7}, {100.4, 131.9}, {101.2, 131.8}, {102.0, 132.0}, {101.8, 131.7}, {101.4, 103.3, 104.7, 105.2, 131.4}, {103.1, 104.1, 105.0, 131.2}, {106.3, 131.5, 132.5}, {107.0, 133.2}, {107.5, 133.7}, {107.8, 133.8}, {107.7, 133.4}, {107.8, 133.2}, {107.8, 133.1}, {107.8, 132.8}, {107.2, 132.5}, {107.0, 132.4}, {107.4, 133.0}, {107.8, 133.9}, {108.1, 134.8}, {108.3, 135.3}, {108.4, 135.2}, {108.2, 135.0}, {108.1, 132.4, 133.3, 135.3}, {108.1, 131.7, 133.0, 134.7}, {108.2, 131.2, 132.7, 134.0}, {108.4, 131.1, 132.9, 133.8}, {108.9, 131.5, 133.2, 134.2}, {109.4, 132.0, 133.7, 134.7}, {109.7, 132.1, 133.8, 134.8}, {109.6, 131.0}, {109.4, 127.7, 128.1, 130.4}, {109.2, 127.3, 128.7, 130.0}, {109.4, 127.5, 129.2, 130.0}, {109.7, 128.1}, {109.0, 128.7}, {109.0, 128.7}, {110.0, 128.1}, {109.6, 111.5, 127.6}, {111.7, 127.8}, {112.3, 128.5}, {113.2, 129.1}, {113.1, 129.2}, {112.7, 129.9}, {112.5, 130.1}, {112.7, 130.5}, {112.9, 130.9}, {112.9, 131.0}, {112.7, 130.9}, {112.7, 130.9}, {113.1, 131.4}, {112.7, 131.8}, {112.4, 131.6}, {113.0, 130.7}, {113.5, 130.1}, {113.2, 129.9}, {113.3, 129.9}, {113.2, 130.4}, {112.4, 131.2}, {113.0, 131.9}, {113.6, 132.6}, {114.1, 132.8}, {114.4, 133.0}, {114.8, 132.9}, {115.2, 132.6}, {116.5, 133.3}, {111.3, 111.9, 116.1, 133.5, 136.2, 136.6}, {109.7, 110.8, 111.6, 115.8, 133.8, 135.7, 136.4}, {109.7, 111.8, 115.8, 134.3, 135.7, 136.6}, {110.2, 112.5, 115.0, 137.3}, {111.0, 113.3, 114.5, 138.4, 140.7}, {111.5, 141.1}, {111.7, 141.2}, {111.9, 141.0}, {112.8, 140.9}, {112.6, 140.7}, {112.7, 114.2, 140.4}, {114.1, 140.5}, {114.1, 140.7, 142.6}, {114.2, 142.8}, {112.7, 114.3, 142.7}, {112.8, 141.3, 142.8}, {112.8, 141.5}, {112.8, 141.5}, {112.7, 141.3}, {112.3, 112.9, 113.6, 141.4}, {112.3, 112.9, 113.9, 141.6}, {112.4, 112.8, 114.1, 141.8}, {114.3, 142.1}, {115.9, 142.5}, {116.1, 143.3}, {116.4, 143.2}, {116.6, 142.8}, {116.5, 141.1}, {116.3, 140.8}, {116.6, 140.9}, {117.1, 141.4}, {117.7, 141.6, 143.9, 144.5}, {118.1, 119.7, 141.5, 143.0, 144.7}, {119.3, 141.5, 142.1, 144.6}, {119.3, 144.8}, {119.7, 145.5}, {118.8, 146.2}, {118.9, 146.4}, {118.4, 146.2}, {118.5, 145.4}, {118.9, 144.5}, {119.0, 144.1}, {119.4, 144.5}, {119.8, 144.8}, {119.7, 144.8}, {118.3, 122.7, 123.3, 144.7}, {117.9, 122.3, 123.4, 126.8, 135.6, 136.2, 144.6}, {118.0, 120.1, 121.6, 127.2, 131.9, 133.3, 135.4, 136.7, 140.0, 144.9}, {118.7, 119.5, 128.1, 129.8, 130.8, 132.3, 134.0, 135.4, 140.7, 145.5}, {129.2, 129.8, 131.9, 132.5, 134.8, 135.5}, {135.5, 135.9}};
		}
	}
}
