netcdf mask {
	:date_created = "20200810T140900";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200810T140900";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 4;
			channels = 1;
			categories = 8;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  15.0, 66.8, 15.0, 60.3;
			max_depth =  72.9,  98.3,  60.3, 115.9;
			start_time = 131315511102200704, 131315511102200704, 131315515112513280, 131315515112513280;
			end_time = 131315515112513280, 131315515112513280, 131315531517357056, 131315531517357056;
			region_id = 1, 2, 3, 4;
			region_name = "Layer1","Layer2","Layer3","Layer4";
			region_provenance = "LSSS", "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "", "";
			region_category_names = "1", "6", "1", "6", "1", "6", "1", "6";
			region_category_proportions = 0.1, 0.9, 0.9, 0.1, 0.1, 0.9, 0.9, 0.1;
			region_category_ids = 1, 2, 3, 4, 5, 6, 7, 8;
			region_type = analysis, analysis, analysis, analysis;
			channel_names = "38";
			region_channels = 1, 1, 1, 1;
			mask_times = {1.313155111022007e+17, 1.313155111125133e+17, 1.313155111228257e+17, 1.313155111332945e+17, 1.31315511143607e+17, 1.313155111539195e+17, 1.313155111647008e+17, 1.313155111747008e+17, 1.313155111851695e+17, 1.313155111956383e+17, 1.31315511206107e+17, 1.313155112165757e+17, 1.313155112270445e+17, 1.313155112372008e+17, 1.313155112473571e+17, 1.313155112582945e+17, 1.313155112690757e+17, 1.313155112795446e+17, 1.31315511289857e+17, 1.313155113006382e+17, 1.313155113106383e+17, 1.313155113211069e+17, 1.313155113325133e+17, 1.313155113431383e+17, 1.313155113540758e+17, 1.313155113642319e+17, 1.313155113748571e+17, 1.313155113851695e+17, 1.313155113953257e+17, 1.313155114056381e+17, 1.313155114157944e+17, 1.313155114264196e+17, 1.313155114364195e+17, 1.313155114564195e+17, 1.313155114673571e+17, 1.313155114781384e+17, 1.313155114882944e+17, 1.313155114989196e+17, 1.313155115095444e+17, 1.313155115200133e+17, 1.313155115311071e+17, 1.313155115412634e+17, 1.313155115515758e+17, 1.31315511561732e+17, 1.313155115718883e+17, 1.313155115822007e+17, 1.31315511592357e+17, 1.313155116031382e+17, 1.313155116140758e+17, 1.313155116247008e+17, 1.313155116348571e+17, 1.313155116451695e+17, 1.31315511655482e+17, 1.31315511666107e+17, 1.313155116772008e+17, 1.313155116873571e+17, 1.313155116981382e+17, 1.313155117090757e+17, 1.31315511719232e+17, 1.313155117297009e+17, 1.31315511739857e+17, 1.313155117509508e+17, 1.31315511761732e+17, 1.313155117718883e+17, 1.313155117820445e+17, 1.313155117926694e+17, 1.313155118037633e+17, 1.313155118140758e+17, 1.313155118243884e+17, 1.313155118345445e+17, 1.31315511845482e+17, 1.313155118556383e+17, 1.313155118664195e+17, 1.313155118772008e+17, 1.313155118876695e+17, 1.313155118982944e+17, 1.313155119095446e+17, 1.313155119206382e+17, 1.313155119307945e+17, 1.313155119409508e+17, 1.313155119518883e+17, 1.313155119625133e+17, 1.313155119731383e+17, 1.313155119831383e+17, 1.31315511993607e+17, 1.313155120039195e+17, 1.313155120140758e+17, 1.313155120250132e+17, 1.313155120353258e+17, 1.313155120457944e+17, 1.313155120568882e+17, 1.313155120670445e+17, 1.313155120776695e+17, 1.313155120882945e+17, 1.313155120984508e+17, 1.313155121089196e+17, 1.31315512119232e+17, 1.313155121297007e+17, 1.313155121403258e+17, 1.313155121507945e+17, 1.313155121612632e+17, 1.31315512172357e+17, 1.31315512182357e+17, 1.313155121928257e+17, 1.31315512202982e+17, 1.313155122142319e+17, 1.313155122248571e+17, 1.313155122350132e+17, 1.313155122456383e+17, 1.313155122559507e+17, 1.31315512266107e+17, 1.313155122762633e+17, 1.313155122864195e+17, 1.313155122964196e+17, 1.313155123075132e+17, 1.313155123178258e+17, 1.313155123284507e+17, 1.31315512339232e+17, 1.313155123497007e+17, 1.313155123597007e+17, 1.31315512370482e+17, 1.313155123806382e+17, 1.313155123909507e+17, 1.313155124018883e+17, 1.313155124122007e+17, 1.313155124226694e+17, 1.313155124332945e+17, 1.31315512443607e+17, 1.313155124540756e+17, 1.313155124642321e+17, 1.31315512474857e+17, 1.313155124853258e+17, 1.31315512495482e+17, 1.313155125057944e+17, 1.31315512516107e+17, 1.313155125265757e+17, 1.313155125373569e+17, 1.313155125482944e+17, 1.31315512559232e+17, 1.313155125693883e+17, 1.313155125797007e+17, 1.313155125903258e+17, 1.313155126006382e+17, 1.313155126206382e+17, 1.313155126309508e+17, 1.313155126412632e+17, 1.313155126515757e+17, 1.313155126618883e+17, 1.313155126722007e+17, 1.313155126828257e+17, 1.313155126937633e+17, 1.313155127039195e+17, 1.313155127140756e+17, 1.313155127242321e+17, 1.313155127343884e+17, 1.313155127447008e+17, 1.31315512755482e+17, 1.313155127659507e+17, 1.313155127762633e+17, 1.313155127864195e+17, 1.313155127965757e+17, 1.31315512806732e+17, 1.313155128170446e+17, 1.313155128272008e+17, 1.313155128372008e+17, 1.313155128475133e+17, 1.313155128584508e+17, 1.313155128697007e+17, 1.313155128803258e+17, 1.313155128906382e+17, 1.313155129011071e+17, 1.31315512911732e+17, 1.31315512922357e+17, 1.313155129326696e+17, 1.313155129428257e+17, 1.313155129534508e+17, 1.31315512963607e+17, 1.313155129743884e+17, 1.313155129845445e+17, 1.31315512995482e+17, 1.313155130062632e+17, 1.313155130164195e+17, 1.31315513026732e+17, 1.313155130368883e+17, 1.313155130472008e+17, 1.313155130573571e+17, 1.313155130681382e+17, 1.313155130782945e+17, 1.313155130887633e+17, 1.31315513099232e+17, 1.31315513109857e+17, 1.31315513120482e+17, 1.313155131312632e+17, 1.313155131420445e+17, 1.313155131525133e+17, 1.313155131634508e+17, 1.313155131739195e+17, 1.313155131842321e+17, 1.313155131945445e+17, 1.313155132047008e+17, 1.313155132153257e+17, 1.313155132259508e+17, 1.31315513236732e+17, 1.313155132484508e+17, 1.313155132589196e+17, 1.313155132703258e+17, 1.313155132806383e+17, 1.313155132906382e+17, 1.313155133026696e+17, 1.313155133134508e+17, 1.31315513323607e+17, 1.313155133343882e+17, 1.313155133450132e+17, 1.313155133556383e+17, 1.313155133657946e+17, 1.313155133762632e+17, 1.313155133865757e+17, 1.313155133972008e+17, 1.313155134076695e+17, 1.313155134182944e+17, 1.313155134284508e+17, 1.31315513439232e+17, 1.313155134493883e+17, 1.313155134593883e+17, 1.31315513469857e+17, 1.313155134801695e+17, 1.313155134903258e+17, 1.313155135006383e+17, 1.313155135115757e+17, 1.313155135225133e+17, 1.313155135331382e+17, 1.313155135432945e+17, 1.31315513553607e+17, 1.313155135637633e+17, 1.313155135742319e+17, 1.313155135842319e+17, 1.313155135951695e+17, 1.313155136062633e+17, 1.31315513616732e+17, 1.313155136273569e+17, 1.313155136378258e+17, 1.313155136482945e+17, 1.31315513658607e+17, 1.313155136690757e+17, 1.313155136797007e+17, 1.313155136901696e+17, 1.313155137009508e+17, 1.313155137112632e+17, 1.313155137215758e+17, 1.313155137318883e+17, 1.313155137426694e+17, 1.313155137528257e+17, 1.313155137632945e+17, 1.313155137742319e+17, 1.313155137845444e+17, 1.313155137947008e+17, 1.313155138048571e+17, 1.31315513815482e+17, 1.313155138257944e+17, 1.313155138364196e+17, 1.313155138465756e+17, 1.313155138568882e+17, 1.313155138668883e+17, 1.313155138778258e+17, 1.313155138882945e+17, 1.313155138987633e+17, 1.31315513909232e+17, 1.313155139200132e+17, 1.313155139303258e+17, 1.313155139407945e+17, 1.313155139512634e+17, 1.313155139615758e+17, 1.313155139720445e+17, 1.313155139826694e+17, 1.313155139931383e+17, 1.313155140034508e+17, 1.313155140136069e+17, 1.313155140243882e+17, 1.313155140353257e+17, 1.313155140468882e+17, 1.313155140573569e+17, 1.313155140675132e+17, 1.313155140781382e+17, 1.313155140884507e+17, 1.313155140990757e+17, 1.313155141092321e+17, 1.31315514119857e+17, 1.313155141300133e+17, 1.313155141500133e+17, 1.313155141601695e+17, 1.313155141703256e+17, 1.313155141806382e+17, 1.313155141907945e+17, 1.313155142009508e+17, 1.313155142112634e+17, 1.313155142215758e+17, 1.31315514232357e+17, 1.313155142426694e+17, 1.31315514252982e+17, 1.313155142632945e+17, 1.313155142834508e+17, 1.313155142937632e+17, 1.313155143040756e+17, 1.313155143147008e+17, 1.313155143251695e+17, 1.313155143359508e+17, 1.31315514346107e+17, 1.313155143562633e+17, 1.313155143670445e+17, 1.313155143775132e+17, 1.313155143884507e+17, 1.313155143987633e+17, 1.313155144089196e+17, 1.313155144193883e+17, 1.313155144301695e+17, 1.313155144403258e+17, 1.313155144504819e+17, 1.313155144618883e+17, 1.313155144722007e+17, 1.313155144832945e+17, 1.313155144936069e+17, 1.313155145043882e+17, 1.313155145147008e+17, 1.313155145251694e+17, 1.31315514535482e+17, 1.313155145456383e+17, 1.313155145557946e+17, 1.313155145659507e+17, 1.313155145762632e+17, 1.313155145870445e+17, 1.313155145982945e+17, 1.313155146087633e+17, 1.313155146195446e+17, 1.31315514629857e+17, 1.313155146401696e+17, 1.31315514650482e+17, 1.313155146606382e+17, 1.313155146717321e+17, 1.31315514681732e+17, 1.31315514692357e+17, 1.313155147025133e+17, 1.313155147126696e+17, 1.313155147231382e+17, 1.313155147337633e+17, 1.313155147442321e+17, 1.313155147547007e+17, 1.313155147651695e+17, 1.313155147753257e+17, 1.313155147856383e+17, 1.313155147959507e+17, 1.313155148073571e+17, 1.313155148182945e+17, 1.313155148287633e+17, 1.313155148397007e+17, 1.31315514850482e+17, 1.31315514860482e+17, 1.313155148714194e+17, 1.313155148818883e+17, 1.313155148931383e+17, 1.313155149034508e+17, 1.313155149139195e+17, 1.313155149243882e+17, 1.313155149348571e+17, 1.313155149451695e+17, 1.313155149557944e+17, 1.313155149659508e+17, 1.31315514976107e+17, 1.313155149868882e+17, 1.313155149972006e+17, 1.313155150075132e+17, 1.313155150178257e+17, 1.313155150279821e+17, 1.313155150390757e+17, 1.313155150497007e+17, 1.313155150603256e+17, 1.31315515070482e+17, 1.313155150809508e+17, 1.313155150915758e+17, 1.313155151018883e+17, 1.313155151125133e+17},
			             {1.313155111022007e+17, 1.313155111125133e+17, 1.313155111228257e+17, 1.313155111332945e+17, 1.31315511143607e+17, 1.313155111539195e+17, 1.313155111647008e+17, 1.313155111747008e+17, 1.313155111851695e+17, 1.313155111956383e+17, 1.31315511206107e+17, 1.313155112165757e+17, 1.313155112270445e+17, 1.313155112372008e+17, 1.313155112473571e+17, 1.313155112582945e+17, 1.313155112690757e+17, 1.313155112795446e+17, 1.31315511289857e+17, 1.313155113006382e+17, 1.313155113106383e+17, 1.313155113211069e+17, 1.313155113325133e+17, 1.313155113431383e+17, 1.313155113540758e+17, 1.313155113642319e+17, 1.313155113748571e+17, 1.313155113851695e+17, 1.313155113953257e+17, 1.313155114056381e+17, 1.313155114157944e+17, 1.313155114264196e+17, 1.313155114364195e+17, 1.313155114564195e+17, 1.313155114673571e+17, 1.313155114781384e+17, 1.313155114882944e+17, 1.313155114989196e+17, 1.313155115095444e+17, 1.313155115200133e+17, 1.313155115311071e+17, 1.313155115412634e+17, 1.313155115515758e+17, 1.31315511561732e+17, 1.313155115718883e+17, 1.313155115822007e+17, 1.31315511592357e+17, 1.313155116031382e+17, 1.313155116140758e+17, 1.313155116247008e+17, 1.313155116348571e+17, 1.313155116451695e+17, 1.31315511655482e+17, 1.31315511666107e+17, 1.313155116772008e+17, 1.313155116873571e+17, 1.313155116981382e+17, 1.313155117090757e+17, 1.31315511719232e+17, 1.313155117297009e+17, 1.31315511739857e+17, 1.313155117509508e+17, 1.31315511761732e+17, 1.313155117718883e+17, 1.313155117820445e+17, 1.313155117926694e+17, 1.313155118037633e+17, 1.313155118140758e+17, 1.313155118243884e+17, 1.313155118345445e+17, 1.31315511845482e+17, 1.313155118556383e+17, 1.313155118664195e+17, 1.313155118772008e+17, 1.313155118876695e+17, 1.313155118982944e+17, 1.313155119095446e+17, 1.313155119206382e+17, 1.313155119307945e+17, 1.313155119409508e+17, 1.313155119518883e+17, 1.313155119625133e+17, 1.313155119731383e+17, 1.313155119831383e+17, 1.31315511993607e+17, 1.313155120039195e+17, 1.313155120140758e+17, 1.313155120250132e+17, 1.313155120353258e+17, 1.313155120457944e+17, 1.313155120568882e+17, 1.313155120670445e+17, 1.313155120776695e+17, 1.313155120882945e+17, 1.313155120984508e+17, 1.313155121089196e+17, 1.31315512119232e+17, 1.313155121297007e+17, 1.313155121403258e+17, 1.313155121507945e+17, 1.313155121612632e+17, 1.31315512172357e+17, 1.31315512182357e+17, 1.313155121928257e+17, 1.31315512202982e+17, 1.313155122142319e+17, 1.313155122248571e+17, 1.313155122350132e+17, 1.313155122456383e+17, 1.313155122559507e+17, 1.31315512266107e+17, 1.313155122762633e+17, 1.313155122864195e+17, 1.313155122964196e+17, 1.313155123075132e+17, 1.313155123178258e+17, 1.313155123284507e+17, 1.31315512339232e+17, 1.313155123497007e+17, 1.313155123597007e+17, 1.31315512370482e+17, 1.313155123806382e+17, 1.313155123909507e+17, 1.313155124018883e+17, 1.313155124122007e+17, 1.313155124226694e+17, 1.313155124332945e+17, 1.31315512443607e+17, 1.313155124540756e+17, 1.313155124642321e+17, 1.31315512474857e+17, 1.313155124853258e+17, 1.31315512495482e+17, 1.313155125057944e+17, 1.31315512516107e+17, 1.313155125265757e+17, 1.313155125373569e+17, 1.313155125482944e+17, 1.31315512559232e+17, 1.313155125693883e+17, 1.313155125797007e+17, 1.313155125903258e+17, 1.313155126006382e+17, 1.313155126206382e+17, 1.313155126309508e+17, 1.313155126412632e+17, 1.313155126515757e+17, 1.313155126618883e+17, 1.313155126722007e+17, 1.313155126828257e+17, 1.313155126937633e+17, 1.313155127039195e+17, 1.313155127140756e+17, 1.313155127242321e+17, 1.313155127343884e+17, 1.313155127447008e+17, 1.31315512755482e+17, 1.313155127659507e+17, 1.313155127762633e+17, 1.313155127864195e+17, 1.313155127965757e+17, 1.31315512806732e+17, 1.313155128170446e+17, 1.313155128272008e+17, 1.313155128372008e+17, 1.313155128475133e+17, 1.313155128584508e+17, 1.313155128697007e+17, 1.313155128803258e+17, 1.313155128906382e+17, 1.313155129011071e+17, 1.31315512911732e+17, 1.31315512922357e+17, 1.313155129326696e+17, 1.313155129428257e+17, 1.313155129534508e+17, 1.31315512963607e+17, 1.313155129743884e+17, 1.313155129845445e+17, 1.31315512995482e+17, 1.313155130062632e+17, 1.313155130164195e+17, 1.31315513026732e+17, 1.313155130368883e+17, 1.313155130472008e+17, 1.313155130573571e+17, 1.313155130681382e+17, 1.313155130782945e+17, 1.313155130887633e+17, 1.31315513099232e+17, 1.31315513109857e+17, 1.31315513120482e+17, 1.313155131312632e+17, 1.313155131420445e+17, 1.313155131525133e+17, 1.313155131634508e+17, 1.313155131739195e+17, 1.313155131842321e+17, 1.313155131945445e+17, 1.313155132047008e+17, 1.313155132153257e+17, 1.313155132259508e+17, 1.31315513236732e+17, 1.313155132484508e+17, 1.313155132589196e+17, 1.313155132703258e+17, 1.313155132806383e+17, 1.313155132906382e+17, 1.313155133026696e+17, 1.313155133134508e+17, 1.31315513323607e+17, 1.313155133343882e+17, 1.313155133450132e+17, 1.313155133556383e+17, 1.313155133657946e+17, 1.313155133762632e+17, 1.313155133865757e+17, 1.313155133972008e+17, 1.313155134076695e+17, 1.313155134182944e+17, 1.313155134284508e+17, 1.31315513439232e+17, 1.313155134493883e+17, 1.313155134593883e+17, 1.31315513469857e+17, 1.313155134801695e+17, 1.313155134903258e+17, 1.313155135006383e+17, 1.313155135115757e+17, 1.313155135225133e+17, 1.313155135331382e+17, 1.313155135432945e+17, 1.31315513553607e+17, 1.313155135637633e+17, 1.313155135742319e+17, 1.313155135842319e+17, 1.313155135951695e+17, 1.313155136062633e+17, 1.31315513616732e+17, 1.313155136273569e+17, 1.313155136378258e+17, 1.313155136482945e+17, 1.31315513658607e+17, 1.313155136690757e+17, 1.313155136797007e+17, 1.313155136901696e+17, 1.313155137009508e+17, 1.313155137112632e+17, 1.313155137215758e+17, 1.313155137318883e+17, 1.313155137426694e+17, 1.313155137528257e+17, 1.313155137632945e+17, 1.313155137742319e+17, 1.313155137845444e+17, 1.313155137947008e+17, 1.313155138048571e+17, 1.31315513815482e+17, 1.313155138257944e+17, 1.313155138364196e+17, 1.313155138465756e+17, 1.313155138568882e+17, 1.313155138668883e+17, 1.313155138778258e+17, 1.313155138882945e+17, 1.313155138987633e+17, 1.31315513909232e+17, 1.313155139200132e+17, 1.313155139303258e+17, 1.313155139407945e+17, 1.313155139512634e+17, 1.313155139615758e+17, 1.313155139720445e+17, 1.313155139826694e+17, 1.313155139931383e+17, 1.313155140034508e+17, 1.313155140136069e+17, 1.313155140243882e+17, 1.313155140353257e+17, 1.313155140468882e+17, 1.313155140573569e+17, 1.313155140675132e+17, 1.313155140781382e+17, 1.313155140884507e+17, 1.313155140990757e+17, 1.313155141092321e+17, 1.31315514119857e+17, 1.313155141300133e+17, 1.313155141500133e+17, 1.313155141601695e+17, 1.313155141703256e+17, 1.313155141806382e+17, 1.313155141907945e+17, 1.313155142009508e+17, 1.313155142112634e+17, 1.313155142215758e+17, 1.31315514232357e+17, 1.313155142426694e+17, 1.31315514252982e+17, 1.313155142632945e+17, 1.313155142834508e+17, 1.313155142937632e+17, 1.313155143040756e+17, 1.313155143147008e+17, 1.313155143251695e+17, 1.313155143359508e+17, 1.31315514346107e+17, 1.313155143562633e+17, 1.313155143670445e+17, 1.313155143775132e+17, 1.313155143884507e+17, 1.313155143987633e+17, 1.313155144089196e+17, 1.313155144193883e+17, 1.313155144301695e+17, 1.313155144403258e+17, 1.313155144504819e+17, 1.313155144618883e+17, 1.313155144722007e+17, 1.313155144832945e+17, 1.313155144936069e+17, 1.313155145043882e+17, 1.313155145147008e+17, 1.313155145251694e+17, 1.31315514535482e+17, 1.313155145456383e+17, 1.313155145557946e+17, 1.313155145659507e+17, 1.313155145762632e+17, 1.313155145870445e+17, 1.313155145982945e+17, 1.313155146087633e+17, 1.313155146195446e+17, 1.31315514629857e+17, 1.313155146401696e+17, 1.31315514650482e+17, 1.313155146606382e+17, 1.313155146717321e+17, 1.31315514681732e+17, 1.31315514692357e+17, 1.313155147025133e+17, 1.313155147126696e+17, 1.313155147231382e+17, 1.313155147337633e+17, 1.313155147442321e+17, 1.313155147547007e+17, 1.313155147651695e+17, 1.313155147753257e+17, 1.313155147856383e+17, 1.313155147959507e+17, 1.313155148073571e+17, 1.313155148182945e+17, 1.313155148287633e+17, 1.313155148397007e+17, 1.31315514850482e+17, 1.31315514860482e+17, 1.313155148714194e+17, 1.313155148818883e+17, 1.313155148931383e+17, 1.313155149034508e+17, 1.313155149139195e+17, 1.313155149243882e+17, 1.313155149348571e+17, 1.313155149451695e+17, 1.313155149557944e+17, 1.313155149659508e+17, 1.31315514976107e+17, 1.313155149868882e+17, 1.313155149972006e+17, 1.313155150075132e+17, 1.313155150178257e+17, 1.313155150279821e+17, 1.313155150390757e+17, 1.313155150497007e+17, 1.313155150603256e+17, 1.31315515070482e+17, 1.313155150809508e+17, 1.313155150915758e+17, 1.313155151018883e+17, 1.313155151125133e+17},
			             {1.313155151125133e+17, 1.313155151226696e+17, 1.31315515132982e+17, 1.313155151434508e+17, 1.313155151550132e+17, 1.313155151653257e+17, 1.31315515175482e+17, 1.313155151857946e+17, 1.313155151959507e+17, 1.313155152065757e+17, 1.313155152175132e+17, 1.31315515227982e+17, 1.313155152382945e+17, 1.313155152487633e+17, 1.313155152593883e+17, 1.313155152700132e+17, 1.313155152807945e+17, 1.313155152911069e+17, 1.313155153022007e+17, 1.313155153126696e+17, 1.313155153232945e+17, 1.313155153334508e+17, 1.313155153439195e+17, 1.313155153542319e+17, 1.31315515364857e+17, 1.313155153751695e+17, 1.313155153856383e+17, 1.313155153957944e+17, 1.31315515406107e+17, 1.313155154173571e+17, 1.313155154281382e+17, 1.313155154390758e+17, 1.313155154501695e+17, 1.31315515460482e+17, 1.31315515471732e+17, 1.313155154825133e+17, 1.313155154926696e+17, 1.313155155032945e+17, 1.313155155134508e+17, 1.313155155240758e+17, 1.31315515534857e+17, 1.313155155451695e+17, 1.313155155559507e+17, 1.313155155665757e+17, 1.313155155765757e+17, 1.313155155875132e+17, 1.313155155976695e+17, 1.313155156078258e+17, 1.313155156184508e+17, 1.313155156293883e+17, 1.313155156397007e+17, 1.313155156501695e+17, 1.313155156607945e+17, 1.313155156714195e+17, 1.313155156818883e+17, 1.313155156928257e+17, 1.31315515702982e+17, 1.313155157131383e+17, 1.31315515723607e+17, 1.313155157340758e+17, 1.313155157442321e+17, 1.313155157543884e+17, 1.313155157651695e+17, 1.313155157757946e+17, 1.31315515786732e+17, 1.313155157968883e+17, 1.313155158072008e+17, 1.313155158173569e+17, 1.313155158275132e+17, 1.313155158376695e+17, 1.313155158479821e+17, 1.31315515857982e+17, 1.313155158681382e+17, 1.313155158789196e+17, 1.313155158890757e+17, 1.313155158995444e+17, 1.313155159103258e+17, 1.313155159211069e+17, 1.313155159312632e+17, 1.313155159414195e+17, 1.31315515952357e+17, 1.313155159625133e+17, 1.31315515972982e+17, 1.31315515982982e+17, 1.313155159931383e+17, 1.313155160039195e+17, 1.31315516014857e+17, 1.313155160251695e+17, 1.31315516035482e+17, 1.31315516046107e+17, 1.313155160565757e+17, 1.313155160668883e+17, 1.313155160776695e+17, 1.313155160881382e+17, 1.313155160984508e+17, 1.313155161086071e+17, 1.31315516119232e+17, 1.31315516129857e+17, 1.313155161411069e+17, 1.313155161522008e+17, 1.313155161625133e+17, 1.313155161728257e+17, 1.313155161831383e+17, 1.313155161937633e+17, 1.313155162039196e+17, 1.313155162143882e+17, 1.313155162247008e+17, 1.313155162356383e+17, 1.313155162462632e+17, 1.31315516256732e+17, 1.313155162668882e+17, 1.313155162772008e+17, 1.313155162875132e+17, 1.313155162978257e+17, 1.313155163081382e+17, 1.313155163182945e+17, 1.313155163284508e+17, 1.31315516339232e+17, 1.313155163501695e+17, 1.313155163603258e+17, 1.313155163706382e+17, 1.313155163811069e+17, 1.313155163912632e+17, 1.313155164014195e+17, 1.313155164115758e+17, 1.313155164215758e+17, 1.313155164326694e+17, 1.313155164428257e+17, 1.313155164531383e+17, 1.313155164639196e+17, 1.313155164745445e+17, 1.313155164847008e+17, 1.313155164953257e+17, 1.313155165062632e+17, 1.313155165164195e+17, 1.313155165270445e+17, 1.313155165375132e+17, 1.313155165478258e+17, 1.313155165581384e+17, 1.313155165684508e+17, 1.313155165787633e+17, 1.31315516589232e+17, 1.313155165993883e+17, 1.313155166097007e+17, 1.313155166200133e+17, 1.31315516630482e+17, 1.313155166409508e+17, 1.313155166514194e+17, 1.313155166615757e+17, 1.313155166718883e+17, 1.313155166831383e+17, 1.31315516693607e+17, 1.313155167045445e+17, 1.313155167150132e+17, 1.313155167253257e+17, 1.313155167362633e+17, 1.313155167462632e+17, 1.313155167564195e+17, 1.313155167675132e+17, 1.313155167784507e+17, 1.31315516788607e+17, 1.313155167989196e+17, 1.31315516809232e+17, 1.313155168195444e+17, 1.313155168297007e+17, 1.313155168403256e+17, 1.31315516850482e+17, 1.313155168612632e+17, 1.313155168714195e+17, 1.313155168820444e+17, 1.313155168922008e+17, 1.313155169037633e+17, 1.313155169143882e+17, 1.313155169245445e+17, 1.313155169351694e+17, 1.31315516945482e+17, 1.313155169568883e+17, 1.313155169672008e+17, 1.313155169776695e+17, 1.313155169887633e+17, 1.31315516999857e+17, 1.313155170101695e+17, 1.31315517020482e+17, 1.313155170307945e+17, 1.313155170411071e+17, 1.313155170514195e+17, 1.313155170618883e+17, 1.313155170720445e+17, 1.313155170822007e+17, 1.313155170931382e+17, 1.313155171037632e+17, 1.313155171139195e+17, 1.313155171242321e+17, 1.313155171343882e+17, 1.313155171447008e+17, 1.313155171551695e+17, 1.31315517166107e+17, 1.313155171765757e+17, 1.313155171868883e+17, 1.313155171970445e+17, 1.313155172170445e+17, 1.313155172278257e+17, 1.313155172382944e+17, 1.313155172484508e+17, 1.313155172589194e+17, 1.313155172693883e+17, 1.313155172795444e+17, 1.313155172900132e+17, 1.313155173006382e+17, 1.313155173109508e+17, 1.313155173214195e+17, 1.313155173315757e+17, 1.313155173418883e+17, 1.31315517352357e+17, 1.313155173626694e+17, 1.31315517372982e+17, 1.313155173832945e+17, 1.31315517393607e+17, 1.313155174039195e+17, 1.313155174142321e+17, 1.313155174243884e+17, 1.313155174347008e+17, 1.31315517444857e+17, 1.313155174551694e+17, 1.313155174653257e+17, 1.313155174757944e+17, 1.313155174865757e+17, 1.313155174978258e+17, 1.313155175082945e+17, 1.313155175193883e+17, 1.31315517529857e+17, 1.31315517540482e+17, 1.313155175507945e+17, 1.31315517562357e+17, 1.313155175725133e+17, 1.313155175837632e+17, 1.313155175940758e+17, 1.313155176042321e+17, 1.313155176143882e+17, 1.313155176243882e+17, 1.313155176345445e+17, 1.313155176453257e+17, 1.31315517656107e+17, 1.313155176665756e+17, 1.313155176768882e+17, 1.313155176872008e+17, 1.313155176973571e+17, 1.31315517707982e+17, 1.313155177184508e+17, 1.313155177290757e+17, 1.313155177395444e+17, 1.31315517749857e+17, 1.313155177600133e+17, 1.313155177704819e+17, 1.313155177807945e+17, 1.313155177912632e+17, 1.313155178017321e+17, 1.313155178122007e+17, 1.31315517822357e+17, 1.313155178325133e+17, 1.31315517842982e+17, 1.313155178534508e+17, 1.313155178639195e+17, 1.313155178747008e+17, 1.313155178850132e+17, 1.313155178959508e+17, 1.31315517906107e+17, 1.313155179165757e+17, 1.313155179273571e+17, 1.313155179375132e+17, 1.313155179482945e+17, 1.31315517958607e+17, 1.313155179687633e+17, 1.313155179793883e+17, 1.313155179895444e+17, 1.31315517999857e+17, 1.31315518009857e+17, 1.313155180200133e+17, 1.313155180307945e+17, 1.313155180411071e+17, 1.313155180514195e+17, 1.313155180617321e+17, 1.313155180718883e+17, 1.313155180822007e+17, 1.31315518092357e+17, 1.313155181028257e+17, 1.31315518112982e+17, 1.313155181232945e+17, 1.313155181340758e+17, 1.313155181442321e+17, 1.313155181543882e+17, 1.313155181645445e+17, 1.313155181753257e+17, 1.31315518185482e+17, 1.313155181957944e+17, 1.313155182065757e+17, 1.313155182172008e+17, 1.313155182273569e+17, 1.31315518237982e+17, 1.31315518247982e+17, 1.313155182584508e+17, 1.313155182695444e+17, 1.313155182801695e+17, 1.313155182904819e+17, 1.313155183012632e+17, 1.313155183115757e+17, 1.31315518322357e+17, 1.313155183325133e+17, 1.313155183428257e+17, 1.313155183531382e+17, 1.313155183634508e+17, 1.313155183747008e+17, 1.31315518386107e+17, 1.31315518396732e+17, 1.313155184075132e+17, 1.31315518417982e+17, 1.313155184284507e+17, 1.31315518438607e+17, 1.313155184492321e+17, 1.313155184595446e+17, 1.31315518469857e+17, 1.313155184801695e+17, 1.313155184907945e+17, 1.313155185014195e+17, 1.313155185122007e+17, 1.313155185226696e+17, 1.313155185326696e+17, 1.313155185439195e+17, 1.313155185545445e+17, 1.313155185645445e+17, 1.31315518575482e+17, 1.313155185856383e+17, 1.313155185959507e+17, 1.31315518606107e+17, 1.313155186173569e+17, 1.313155186276695e+17, 1.313155186378257e+17, 1.31315518648607e+17, 1.313155186595446e+17, 1.313155186701695e+17, 1.313155186806383e+17, 1.313155186909508e+17, 1.313155187011069e+17, 1.313155187115757e+17, 1.31315518721732e+17, 1.313155187318883e+17, 1.31315518742357e+17, 1.313155187525133e+17, 1.313155187628257e+17, 1.313155187739195e+17, 1.313155187840758e+17, 1.313155187945445e+17, 1.313155188047008e+17, 1.313155188150132e+17, 1.313155188253258e+17, 1.31315518836732e+17, 1.313155188476695e+17, 1.313155188578257e+17, 1.31315518867982e+17, 1.313155188782945e+17, 1.313155188884508e+17, 1.313155188987633e+17, 1.313155189090757e+17, 1.313155189195446e+17, 1.313155189303258e+17, 1.31315518940482e+17, 1.313155189506383e+17, 1.313155189607945e+17, 1.313155189714195e+17, 1.313155189815758e+17, 1.313155189918883e+17, 1.31315519002357e+17, 1.313155190126696e+17, 1.313155190232946e+17, 1.31315519033607e+17, 1.313155190439195e+17, 1.313155190542321e+17, 1.31315519064857e+17, 1.313155190750132e+17, 1.313155190850132e+17, 1.313155190953257e+17, 1.313155191059508e+17, 1.31315519116107e+17, 1.313155191264195e+17, 1.313155191365757e+17, 1.31315519146732e+17, 1.313155191570445e+17, 1.313155191681382e+17, 1.313155191784508e+17, 1.313155191887633e+17, 1.313155191987633e+17, 1.313155192089196e+17, 1.313155192195446e+17, 1.31315519229857e+17, 1.31315519240482e+17, 1.313155192506383e+17, 1.313155192612632e+17, 1.313155192714195e+17, 1.31315519281732e+17, 1.313155192920444e+17, 1.313155193026694e+17, 1.313155193126696e+17, 1.31315519323607e+17, 1.313155193340758e+17, 1.313155193445444e+17, 1.313155193550132e+17, 1.31315519365482e+17, 1.313155193757946e+17, 1.31315519386107e+17, 1.313155193964196e+17, 1.31315519406732e+17, 1.313155194168882e+17, 1.313155194273571e+17, 1.313155194376695e+17, 1.313155194484507e+17, 1.313155194590757e+17, 1.31315519469232e+17, 1.313155194800132e+17, 1.313155194901695e+17, 1.31315519500482e+17, 1.313155195106383e+17, 1.313155195211069e+17, 1.31315519531732e+17, 1.313155195418883e+17, 1.31315519552357e+17, 1.313155195625133e+17, 1.313155195726696e+17, 1.313155195832945e+17, 1.313155195940758e+17, 1.31315519605482e+17, 1.313155196157944e+17, 1.31315519626107e+17, 1.313155196372008e+17, 1.313155196476695e+17, 1.31315519657982e+17, 1.313155196681382e+17, 1.31315519678607e+17, 1.313155196889196e+17, 1.313155196989196e+17, 1.313155197093883e+17, 1.313155197203258e+17, 1.31315519730482e+17, 1.313155197409508e+17, 1.313155197512632e+17, 1.31315519761732e+17, 1.313155197720444e+17, 1.313155197825133e+17, 1.313155197926696e+17, 1.313155198032945e+17, 1.313155198140758e+17, 1.313155198242321e+17, 1.313155198345445e+17, 1.313155198450132e+17, 1.31315519855482e+17, 1.31315519866107e+17, 1.31315519876732e+17, 1.313155198878258e+17, 1.313155198984507e+17, 1.313155199089194e+17, 1.313155199195446e+17, 1.313155199306382e+17, 1.313155199420445e+17, 1.313155199522008e+17, 1.31315519962357e+17, 1.313155199726694e+17, 1.313155199828257e+17, 1.31315519992982e+17, 1.313155200037632e+17, 1.313155200150132e+17, 1.313155200251695e+17, 1.313155200353257e+17, 1.313155200456383e+17, 1.313155200562633e+17, 1.313155200664196e+17, 1.313155200772006e+17, 1.31315520087982e+17, 1.31315520098607e+17, 1.31315520109232e+17, 1.313155201193883e+17, 1.313155201297007e+17, 1.31315520140482e+17, 1.313155201506382e+17, 1.313155201607945e+17, 1.313155201714195e+17, 1.313155201822007e+17, 1.313155201925133e+17, 1.313155202026696e+17, 1.313155202134508e+17, 1.313155202236069e+17, 1.313155202337632e+17, 1.313155202439195e+17, 1.313155202550132e+17, 1.313155202653257e+17, 1.313155202754821e+17, 1.313155202868883e+17, 1.313155202972008e+17, 1.313155203073569e+17, 1.313155203178258e+17, 1.313155203282945e+17, 1.31315520339232e+17, 1.313155203495444e+17, 1.31315520359857e+17, 1.313155203704819e+17, 1.313155203811071e+17, 1.313155203914195e+17, 1.313155204014195e+17, 1.313155204115757e+17, 1.313155204225133e+17, 1.313155204326696e+17, 1.313155204437633e+17, 1.313155204540758e+17, 1.313155204643884e+17, 1.313155204750132e+17, 1.313155204850132e+17, 1.313155204953258e+17, 1.313155205057944e+17, 1.313155205162633e+17, 1.313155205264196e+17, 1.313155205365757e+17, 1.313155205468883e+17, 1.313155205570445e+17, 1.313155205676695e+17, 1.313155205789196e+17, 1.313155205900133e+17, 1.31315520600482e+17, 1.313155206112632e+17, 1.313155206215757e+17, 1.313155206318883e+17, 1.313155206422007e+17, 1.313155206526696e+17, 1.31315520663607e+17, 1.313155206743882e+17, 1.313155206847007e+17, 1.313155206951695e+17, 1.313155207057944e+17, 1.313155207165757e+17, 1.313155207270445e+17, 1.31315520737982e+17, 1.31315520748607e+17, 1.313155207587633e+17, 1.313155207689196e+17, 1.313155207793882e+17, 1.313155207900133e+17, 1.313155208007945e+17, 1.313155208112634e+17, 1.31315520821732e+17, 1.313155208326696e+17, 1.31315520842982e+17, 1.31315520852982e+17, 1.313155208634508e+17, 1.313155208740756e+17, 1.313155208842321e+17, 1.313155208943882e+17, 1.313155209047008e+17, 1.313155209150132e+17, 1.313155209253257e+17, 1.31315520936107e+17, 1.31315520946732e+17, 1.313155209575132e+17, 1.313155209675133e+17, 1.313155209781382e+17, 1.31315520988607e+17, 1.313155209997007e+17, 1.313155210107945e+17, 1.313155210211069e+17, 1.313155210311071e+17, 1.313155210412632e+17, 1.313155210514195e+17, 1.31315521061732e+17, 1.31315521072357e+17, 1.313155210826694e+17, 1.31315521092982e+17, 1.313155211037632e+17, 1.313155211140758e+17, 1.313155211248571e+17, 1.31315521136107e+17, 1.31315521146732e+17, 1.313155211568883e+17, 1.313155211672008e+17, 1.313155211773569e+17, 1.313155211878258e+17, 1.313155211982945e+17, 1.313155212087633e+17, 1.313155212200133e+17, 1.31315521230482e+17, 1.313155212407945e+17, 1.313155212511071e+17, 1.313155212622007e+17, 1.313155212725133e+17, 1.313155212839196e+17, 1.313155212943882e+17, 1.31315521304857e+17, 1.313155213153257e+17, 1.31315521325482e+17, 1.313155213357944e+17, 1.31315521346107e+17, 1.31315521356732e+17, 1.313155213678258e+17, 1.313155213781382e+17, 1.313155213884508e+17, 1.31315521398607e+17, 1.313155214087633e+17, 1.313155214287633e+17, 1.313155214393883e+17, 1.313155214500132e+17, 1.313155214609508e+17, 1.313155214712632e+17, 1.313155214815757e+17, 1.313155214918883e+17, 1.313155215022007e+17, 1.31315521512357e+17, 1.313155215226696e+17, 1.31315521533607e+17, 1.313155215439196e+17, 1.313155215547007e+17, 1.31315521564857e+17, 1.313155215764195e+17, 1.31315521586732e+17, 1.313155215976695e+17, 1.31315521607982e+17, 1.313155216182945e+17, 1.313155216287631e+17, 1.313155216389194e+17, 1.31315521649232e+17, 1.313155216595444e+17, 1.313155216700132e+17, 1.313155216807945e+17, 1.313155216912632e+17, 1.313155217012634e+17, 1.313155217115758e+17, 1.313155217218883e+17, 1.313155217325133e+17, 1.313155217434508e+17, 1.31315521753607e+17, 1.31315521764857e+17, 1.313155217750132e+17, 1.313155217851695e+17, 1.313155217953258e+17, 1.31315521805482e+17, 1.313155218159507e+17, 1.31315521826107e+17, 1.313155218362633e+17, 1.313155218465757e+17, 1.313155218578257e+17, 1.313155218682945e+17, 1.313155218789196e+17, 1.313155218897007e+17, 1.31315521899857e+17, 1.313155219101696e+17, 1.313155219212632e+17, 1.313155219315757e+17, 1.313155219418883e+17, 1.31315521952357e+17, 1.313155219626694e+17, 1.313155219737632e+17, 1.313155219839195e+17, 1.313155219939195e+17, 1.313155220040758e+17, 1.313155220143882e+17, 1.313155220250134e+17, 1.313155220351695e+17, 1.313155220453257e+17, 1.313155220556383e+17, 1.31315522066107e+17, 1.313155220764195e+17, 1.313155220867319e+17, 1.313155220968882e+17, 1.313155221075132e+17, 1.313155221182944e+17, 1.313155221293883e+17, 1.313155221401695e+17, 1.313155221509508e+17, 1.313155221611071e+17, 1.31315522171732e+17, 1.313155221828257e+17, 1.31315522192982e+17, 1.313155222039195e+17, 1.313155222140758e+17, 1.313155222245445e+17, 1.313155222353258e+17, 1.313155222464195e+17, 1.31315522256732e+17, 1.313155222672006e+17, 1.313155222773569e+17, 1.313155222875132e+17, 1.313155222989196e+17, 1.313155223097007e+17, 1.31315522319857e+17, 1.313155223303256e+17, 1.31315522340482e+17, 1.313155223511069e+17, 1.313155223612632e+17, 1.313155223714195e+17, 1.313155223820444e+17, 1.313155223920445e+17, 1.31315522402982e+17, 1.31315522413607e+17, 1.313155224237633e+17, 1.313155224342319e+17, 1.313155224442321e+17, 1.31315522454857e+17, 1.313155224650132e+17, 1.313155224751695e+17, 1.31315522485482e+17, 1.313155224957946e+17, 1.31315522506107e+17, 1.313155225162633e+17, 1.313155225264196e+17, 1.31315522536732e+17, 1.313155225470445e+17, 1.313155225578258e+17, 1.313155225682945e+17, 1.313155225784508e+17, 1.313155225887633e+17, 1.313155225993883e+17, 1.313155226104819e+17, 1.313155226214194e+17, 1.31315522631732e+17, 1.313155226420444e+17, 1.31315522652357e+17, 1.313155226628257e+17, 1.313155226742319e+17, 1.313155226843882e+17, 1.313155226945445e+17, 1.313155227047007e+17, 1.31315522714857e+17, 1.313155227253257e+17, 1.313155227359507e+17, 1.313155227462633e+17, 1.313155227564196e+17, 1.313155227668883e+17, 1.313155227773571e+17, 1.313155227876695e+17, 1.313155227984508e+17, 1.31315522808607e+17, 1.313155228193882e+17, 1.313155228295444e+17, 1.31315522839857e+17, 1.313155228503258e+17, 1.313155228612632e+17, 1.313155228726696e+17, 1.313155228831382e+17, 1.313155228934508e+17, 1.313155229045445e+17, 1.313155229151695e+17, 1.313155229262633e+17, 1.313155229365757e+17, 1.31315522947982e+17, 1.313155229584508e+17, 1.313155229690758e+17, 1.313155229804819e+17, 1.313155229911071e+17, 1.313155230022007e+17, 1.31315523012357e+17, 1.313155230228257e+17, 1.31315523032982e+17, 1.313155230431383e+17, 1.313155230534508e+17, 1.313155230642319e+17, 1.313155230743882e+17, 1.313155230847008e+17, 1.313155230953257e+17, 1.31315523105482e+17, 1.313155231156383e+17, 1.313155231270445e+17, 1.313155231379821e+17, 1.313155231484508e+17, 1.313155231592321e+17, 1.31315523169857e+17, 1.313155231801695e+17, 1.313155231906382e+17, 1.313155232011071e+17, 1.313155232114195e+17, 1.313155232214195e+17, 1.313155232318883e+17, 1.313155232418883e+17, 1.313155232525133e+17, 1.313155232634508e+17, 1.313155232739195e+17, 1.313155232842319e+17, 1.313155232945445e+17, 1.31315523304857e+17, 1.313155233150132e+17, 1.313155233251695e+17, 1.313155233353257e+17, 1.31315523345482e+17, 1.313155233556383e+17, 1.31315523366107e+17, 1.313155233764195e+17, 1.313155233865757e+17, 1.313155233973571e+17, 1.313155234078258e+17, 1.313155234179821e+17, 1.31315523428607e+17, 1.313155234390757e+17, 1.31315523449232e+17, 1.31315523459232e+17, 1.31315523469857e+17, 1.313155234800133e+17, 1.313155234911069e+17, 1.313155235014195e+17, 1.313155235126694e+17, 1.313155235236069e+17, 1.313155235343882e+17, 1.31315523544857e+17, 1.313155235556383e+17, 1.313155235657946e+17, 1.313155235765757e+17, 1.313155235870445e+17, 1.313155235975132e+17, 1.313155236081382e+17, 1.31315523618607e+17, 1.313155236289196e+17, 1.31315523639232e+17, 1.313155236593883e+17, 1.313155236695446e+17, 1.313155236797007e+17, 1.313155236900132e+17, 1.313155237003256e+17, 1.313155237106382e+17, 1.313155237209508e+17, 1.313155237309508e+17, 1.313155237414195e+17, 1.313155237515758e+17, 1.313155237618883e+17, 1.313155237720444e+17, 1.313155237825133e+17, 1.313155237928257e+17, 1.313155238037633e+17, 1.313155238142321e+17, 1.313155238243882e+17, 1.313155238345444e+17, 1.313155238447008e+17, 1.313155238548571e+17, 1.313155238653257e+17, 1.313155238765757e+17, 1.31315523886732e+17, 1.313155238976695e+17, 1.313155239078258e+17, 1.313155239187633e+17, 1.313155239297007e+17, 1.313155239400133e+17, 1.313155239514195e+17, 1.313155239615757e+17, 1.313155239725133e+17, 1.31315523982982e+17, 1.313155239934508e+17, 1.313155240037633e+17, 1.313155240142321e+17, 1.31315524025482e+17, 1.313155240359507e+17, 1.313155240462633e+17, 1.313155240570445e+17, 1.313155240675132e+17, 1.31315524078607e+17, 1.31315524089232e+17, 1.31315524099232e+17, 1.313155241095444e+17, 1.31315524119857e+17, 1.313155241301695e+17, 1.313155241406382e+17, 1.313155241507945e+17, 1.313155241609508e+17, 1.313155241714195e+17, 1.313155241815758e+17, 1.313155241926696e+17, 1.313155242032945e+17, 1.313155242134508e+17, 1.313155242242321e+17, 1.313155242345445e+17, 1.313155242450132e+17, 1.313155242551695e+17, 1.313155242657944e+17, 1.31315524276732e+17, 1.313155242870445e+17, 1.313155242978258e+17, 1.313155243090757e+17, 1.313155243193883e+17, 1.313155243301695e+17, 1.313155243406382e+17, 1.313155243514195e+17, 1.313155243615758e+17, 1.313155243715757e+17, 1.313155243818883e+17, 1.313155243922007e+17, 1.313155244025133e+17, 1.313155244139195e+17, 1.313155244240758e+17, 1.31315524434857e+17, 1.313155244451695e+17, 1.313155244553257e+17, 1.313155244656383e+17, 1.31315524476107e+17, 1.313155244862633e+17, 1.313155244973569e+17, 1.313155245082944e+17, 1.313155245184508e+17, 1.313155245286071e+17, 1.313155245395444e+17, 1.313155245501695e+17, 1.313155245609508e+17, 1.313155245718883e+17, 1.31315524582357e+17, 1.313155245928257e+17, 1.313155246032945e+17, 1.313155246134508e+17, 1.31315524623607e+17, 1.313155246340756e+17, 1.313155246442321e+17, 1.313155246543884e+17, 1.313155246647008e+17, 1.313155246750132e+17, 1.313155246857944e+17, 1.31315524696107e+17, 1.31315524706732e+17, 1.313155247168883e+17, 1.313155247281382e+17, 1.31315524738607e+17, 1.313155247489194e+17, 1.313155247603258e+17, 1.313155247711071e+17, 1.31315524781732e+17, 1.313155247922008e+17, 1.313155248028257e+17, 1.31315524813607e+17, 1.313155248239195e+17, 1.313155248340758e+17, 1.313155248445445e+17, 1.31315524855482e+17, 1.313155248657946e+17, 1.313155248762633e+17, 1.313155248870445e+17, 1.313155248973571e+17, 1.313155249075132e+17, 1.313155249178257e+17, 1.313155249282945e+17, 1.313155249392321e+17, 1.313155249493883e+17, 1.31315524959857e+17, 1.313155249700132e+17, 1.313155249803258e+17, 1.313155249912632e+17, 1.313155250022007e+17, 1.313155250126696e+17, 1.313155250232945e+17, 1.31315525033607e+17, 1.313155250437633e+17, 1.313155250543882e+17, 1.313155250645445e+17, 1.31315525074857e+17, 1.31315525085482e+17, 1.313155250962632e+17, 1.313155251064195e+17, 1.313155251165757e+17, 1.313155251265757e+17, 1.313155251370445e+17, 1.313155251476695e+17, 1.313155251586071e+17, 1.313155251690757e+17, 1.31315525179232e+17, 1.313155251893882e+17, 1.313155251997007e+17, 1.313155252100132e+17, 1.313155252201695e+17, 1.313155252311069e+17, 1.313155252415757e+17, 1.313155252520445e+17, 1.31315525262357e+17, 1.313155252734508e+17, 1.313155252843884e+17, 1.313155252947008e+17, 1.31315525304857e+17, 1.313155253153258e+17, 1.313155253259507e+17, 1.31315525336732e+17, 1.313155253470445e+17, 1.313155253572008e+17, 1.313155253676695e+17, 1.313155253784508e+17, 1.31315525388607e+17, 1.313155254001695e+17, 1.313155254106383e+17, 1.313155254206382e+17, 1.313155254311069e+17, 1.313155254414194e+17, 1.313155254518883e+17, 1.31315525462357e+17, 1.313155254726696e+17, 1.313155254831383e+17, 1.313155254934508e+17, 1.313155255037633e+17, 1.313155255142319e+17, 1.313155255243882e+17, 1.313155255345445e+17, 1.31315525545482e+17, 1.313155255559507e+17, 1.313155255664195e+17, 1.31315525576732e+17, 1.313155255868883e+17, 1.313155255970445e+17, 1.313155256073569e+17, 1.313155256176695e+17, 1.313155256278258e+17, 1.313155256382944e+17, 1.313155256484507e+17, 1.31315525658607e+17, 1.313155256693883e+17, 1.31315525679857e+17, 1.313155256900133e+17, 1.313155257006383e+17, 1.313155257109508e+17, 1.313155257212632e+17, 1.313155257314195e+17, 1.313155257417321e+17, 1.31315525752357e+17, 1.313155257628257e+17, 1.313155257734508e+17, 1.313155257842321e+17, 1.313155257951695e+17, 1.313155258053257e+17, 1.31315525815482e+17, 1.313155258257946e+17, 1.313155258370445e+17, 1.313155258475132e+17, 1.313155258579821e+17, 1.313155258682945e+17, 1.31315525879232e+17, 1.31315525889857e+17, 1.313155259003258e+17, 1.313155259103258e+17, 1.313155259206382e+17, 1.313155259311069e+17, 1.313155259412632e+17, 1.31315525952357e+17, 1.313155259632945e+17, 1.31315525973607e+17, 1.313155259837633e+17, 1.313155259942319e+17, 1.313155260043882e+17, 1.313155260145445e+17, 1.313155260250132e+17, 1.313155260353257e+17, 1.313155260457944e+17, 1.31315526056107e+17, 1.313155260665757e+17, 1.313155260773571e+17, 1.313155260875133e+17, 1.313155260982945e+17, 1.313155261095444e+17, 1.31315526119857e+17, 1.31315526130482e+17, 1.313155261407945e+17, 1.313155261509507e+17, 1.313155261611069e+17, 1.313155261714195e+17, 1.313155261825133e+17, 1.31315526192982e+17, 1.313155262031383e+17, 1.313155262134508e+17, 1.313155262240758e+17, 1.313155262359507e+17, 1.31315526246107e+17, 1.313155262564195e+17, 1.31315526266732e+17, 1.31315526277982e+17, 1.313155262882944e+17, 1.31315526298607e+17, 1.31315526309232e+17, 1.313155263193883e+17, 1.313155263297007e+17, 1.313155263400132e+17, 1.313155263506382e+17, 1.313155263611069e+17, 1.313155263712632e+17, 1.313155263815757e+17, 1.313155263926696e+17, 1.31315526402982e+17, 1.313155264132945e+17, 1.31315526423607e+17, 1.313155264337633e+17, 1.313155264445445e+17, 1.31315526454857e+17, 1.313155264657946e+17, 1.31315526476107e+17, 1.313155264864195e+17, 1.313155264970445e+17, 1.313155265073571e+17, 1.313155265181382e+17, 1.313155265287633e+17, 1.313155265395444e+17, 1.313155265509508e+17, 1.313155265611069e+17, 1.313155265715758e+17, 1.313155265822007e+17, 1.313155265925133e+17, 1.313155266037633e+17, 1.313155266140758e+17, 1.313155266243882e+17, 1.313155266347008e+17, 1.31315526644857e+17, 1.313155266553257e+17, 1.313155266659507e+17, 1.31315526676107e+17, 1.313155266864196e+17, 1.313155266973571e+17, 1.313155267078258e+17, 1.313155267184507e+17, 1.313155267290757e+17, 1.31315526740482e+17, 1.313155267507945e+17, 1.313155267618883e+17, 1.313155267720445e+17, 1.31315526782357e+17, 1.313155267925133e+17, 1.313155268032945e+17, 1.31315526813607e+17, 1.313155268237633e+17, 1.313155268339195e+17, 1.313155268442319e+17, 1.31315526855482e+17, 1.313155268672008e+17, 1.31315526877982e+17, 1.31315526888607e+17, 1.31315526899232e+17, 1.313155269093883e+17, 1.31315526919857e+17, 1.313155269301696e+17, 1.31315526940482e+17, 1.313155269507945e+17, 1.313155269609508e+17, 1.313155269712632e+17, 1.31315526982982e+17, 1.313155269936069e+17, 1.313155270045445e+17, 1.31315527014857e+17, 1.313155270257944e+17, 1.313155270359507e+17, 1.313155270462633e+17, 1.313155270565757e+17, 1.313155270673571e+17, 1.313155270778258e+17, 1.313155270882944e+17, 1.31315527098607e+17, 1.313155271087633e+17, 1.31315527119232e+17, 1.313155271295444e+17, 1.313155271400132e+17, 1.313155271506383e+17, 1.313155271614195e+17, 1.313155271715757e+17, 1.313155271822008e+17, 1.31315527193607e+17, 1.313155272042321e+17, 1.313155272147007e+17, 1.313155272250132e+17, 1.313155272353257e+17, 1.31315527245482e+17, 1.313155272557944e+17, 1.31315527266107e+17, 1.313155272764196e+17, 1.313155272873571e+17, 1.313155272976695e+17, 1.313155273082944e+17, 1.313155273184507e+17, 1.313155273290757e+17, 1.313155273395446e+17, 1.313155273501695e+17, 1.313155273603258e+17, 1.313155273706383e+17, 1.313155273809508e+17, 1.313155273911071e+17, 1.31315527401732e+17, 1.31315527412357e+17, 1.313155274225133e+17, 1.313155274331383e+17, 1.313155274431382e+17, 1.313155274540758e+17, 1.313155274642321e+17, 1.313155274745445e+17, 1.313155274845445e+17, 1.313155274959507e+17, 1.31315527506107e+17, 1.313155275162633e+17, 1.313155275265757e+17, 1.313155275367319e+17, 1.313155275472008e+17, 1.313155275575132e+17, 1.313155275679821e+17, 1.313155275782945e+17, 1.313155275897007e+17, 1.313155276003258e+17, 1.313155276114195e+17, 1.31315527622357e+17, 1.313155276323571e+17, 1.31315527643607e+17, 1.313155276539195e+17, 1.313155276642319e+17, 1.313155276745445e+17, 1.313155276851695e+17, 1.31315527696107e+17, 1.313155277062632e+17, 1.313155277165757e+17, 1.31315527726732e+17, 1.313155277368883e+17, 1.313155277476695e+17, 1.31315527758607e+17, 1.313155277690757e+17, 1.313155277800133e+17, 1.313155277903258e+17, 1.31315527801732e+17, 1.313155278126696e+17, 1.313155278237633e+17, 1.313155278340758e+17, 1.313155278450132e+17, 1.31315527856107e+17, 1.31315527866732e+17, 1.313155278778258e+17, 1.313155278884507e+17, 1.313155278989196e+17, 1.313155279093883e+17, 1.313155279195444e+17, 1.313155279301695e+17, 1.313155279403258e+17, 1.313155279509508e+17, 1.313155279609508e+17, 1.313155279718883e+17, 1.313155279820444e+17, 1.313155279922007e+17, 1.31315528002357e+17, 1.313155280125133e+17, 1.313155280237633e+17, 1.313155280339196e+17, 1.313155280440758e+17, 1.31315528054857e+17, 1.313155280654821e+17, 1.313155280759507e+17, 1.313155280862633e+17, 1.313155280972008e+17, 1.313155281075132e+17, 1.313155281178258e+17, 1.313155281279821e+17, 1.313155281382945e+17, 1.313155281495444e+17, 1.313155281600132e+17, 1.313155281703258e+17, 1.313155281807945e+17, 1.313155281911069e+17, 1.313155282012632e+17, 1.313155282128257e+17, 1.313155282242319e+17, 1.313155282345445e+17, 1.313155282456383e+17, 1.313155282562633e+17, 1.313155282664195e+17, 1.313155282765757e+17, 1.31315528286732e+17, 1.313155282975133e+17, 1.313155283082944e+17, 1.31315528318607e+17, 1.313155283287633e+17, 1.313155283389196e+17, 1.313155283495444e+17, 1.313155283607945e+17, 1.313155283709508e+17, 1.313155283814195e+17, 1.313155283931383e+17, 1.313155284034508e+17, 1.31315528413607e+17, 1.313155284239195e+17, 1.313155284343882e+17, 1.313155284445445e+17, 1.313155284553257e+17, 1.313155284662632e+17, 1.313155284764195e+17, 1.313155284868882e+17, 1.313155284972006e+17, 1.313155285075132e+17, 1.313155285182945e+17, 1.313155285290757e+17, 1.313155285395444e+17, 1.31315528549857e+17, 1.31315528559857e+17, 1.313155285701695e+17, 1.313155285803258e+17, 1.313155285907945e+17, 1.313155286020444e+17, 1.31315528612357e+17, 1.313155286232945e+17, 1.313155286342321e+17, 1.31315528645482e+17, 1.313155286557944e+17, 1.313155286657944e+17, 1.313155286765757e+17, 1.313155286868883e+17, 1.313155286970445e+17, 1.31315528707982e+17, 1.313155287193883e+17, 1.313155287301695e+17, 1.313155287407944e+17, 1.313155287512632e+17, 1.313155287618883e+17, 1.313155287720445e+17, 1.313155287825133e+17, 1.313155287932945e+17, 1.31315528803607e+17, 1.313155288137632e+17, 1.313155288247007e+17, 1.313155288357946e+17, 1.313155288462633e+17, 1.313155288570445e+17, 1.313155288675133e+17, 1.313155288784508e+17, 1.313155288889196e+17, 1.31315528899857e+17, 1.313155289115757e+17, 1.31315528921732e+17, 1.313155289318883e+17, 1.313155289431382e+17, 1.313155289534508e+17, 1.313155289637632e+17, 1.313155289740756e+17, 1.313155289842321e+17, 1.313155289945445e+17, 1.31315529004857e+17, 1.313155290153257e+17, 1.313155290253258e+17, 1.31315529035482e+17, 1.313155290457944e+17, 1.313155290572008e+17, 1.313155290676695e+17, 1.313155290778258e+17, 1.313155290879821e+17, 1.313155290982945e+17, 1.313155291084507e+17, 1.313155291193883e+17, 1.313155291295444e+17, 1.31315529139857e+17, 1.31315529150482e+17, 1.313155291612632e+17, 1.313155291715757e+17, 1.31315529181732e+17, 1.313155291922007e+17, 1.313155292028257e+17, 1.313155292142321e+17, 1.313155292251695e+17, 1.313155292362633e+17, 1.313155292464196e+17, 1.313155292565757e+17, 1.313155292670445e+17, 1.313155292773571e+17, 1.313155292875132e+17, 1.31315529297982e+17, 1.313155293079821e+17, 1.313155293182945e+17, 1.313155293290757e+17, 1.313155293401695e+17, 1.313155293511069e+17, 1.313155293612632e+17, 1.313155293714194e+17, 1.313155293818883e+17, 1.313155293922008e+17, 1.31315529402357e+17, 1.313155294125133e+17, 1.313155294226696e+17, 1.313155294331383e+17, 1.313155294434508e+17, 1.313155294543882e+17, 1.313155294651695e+17, 1.313155294765757e+17, 1.31315529487982e+17, 1.313155294981382e+17, 1.313155295084507e+17, 1.313155295187633e+17, 1.313155295287631e+17, 1.313155295393883e+17, 1.313155295495446e+17, 1.31315529559857e+17, 1.313155295700132e+17, 1.313155295801695e+17, 1.313155295907945e+17, 1.313155296012634e+17, 1.313155296115758e+17, 1.313155296225133e+17, 1.31315529632982e+17, 1.313155296434508e+17, 1.313155296540758e+17, 1.313155296651695e+17, 1.313155296751695e+17, 1.313155296853257e+17, 1.313155296956383e+17, 1.313155297056383e+17, 1.313155297159507e+17, 1.313155297265757e+17, 1.31315529736732e+17, 1.313155297482945e+17, 1.313155297593883e+17, 1.31315529769857e+17, 1.313155297803258e+17, 1.313155297911069e+17, 1.313155298012632e+17, 1.313155298118883e+17, 1.313155298220444e+17, 1.313155298326696e+17, 1.313155298437633e+17, 1.313155298539195e+17, 1.313155298642321e+17, 1.313155298743882e+17, 1.313155298847007e+17, 1.313155298953257e+17, 1.313155299057946e+17, 1.313155299159508e+17, 1.31315529926107e+17, 1.313155299362633e+17, 1.313155299464196e+17, 1.313155299565757e+17, 1.31315529966732e+17, 1.313155299775132e+17, 1.313155299878257e+17, 1.313155299981382e+17, 1.313155300090757e+17, 1.31315530019857e+17, 1.313155300301695e+17, 1.313155300403258e+17, 1.313155300507945e+17, 1.313155300614195e+17, 1.313155300722008e+17, 1.313155300823571e+17, 1.313155300928257e+17, 1.31315530102982e+17, 1.313155301131382e+17, 1.313155301232945e+17, 1.313155301340758e+17, 1.313155301457944e+17, 1.313155301564195e+17, 1.31315530166732e+17, 1.313155301768882e+17, 1.313155301872008e+17, 1.313155301976695e+17, 1.313155302078257e+17, 1.313155302182944e+17, 1.313155302284508e+17, 1.313155302397009e+17, 1.313155302500133e+17, 1.313155302603258e+17, 1.313155302704819e+17, 1.313155302812632e+17, 1.313155302920445e+17, 1.31315530302357e+17, 1.313155303126696e+17, 1.31315530322982e+17, 1.313155303331382e+17, 1.313155303437632e+17, 1.313155303539195e+17, 1.313155303640756e+17, 1.313155303743882e+17, 1.313155303845445e+17, 1.313155303947008e+17, 1.313155304056383e+17, 1.313155304159507e+17, 1.313155304265757e+17, 1.313155304368882e+17, 1.313155304472008e+17, 1.313155304575132e+17, 1.313155304687633e+17, 1.313155304789194e+17, 1.31315530489232e+17, 1.313155304997007e+17, 1.313155305104819e+17, 1.31315530520482e+17, 1.313155305306382e+17, 1.313155305407945e+17, 1.313155305514195e+17, 1.313155305617321e+17, 1.313155305720445e+17, 1.313155305822007e+17, 1.31315530592357e+17, 1.313155306025133e+17, 1.313155306128257e+17, 1.31315530622982e+17, 1.313155306331382e+17, 1.313155306440758e+17, 1.313155306543882e+17, 1.313155306659507e+17, 1.313155306765757e+17, 1.31315530686732e+17, 1.313155306972008e+17, 1.313155307075133e+17, 1.313155307181382e+17, 1.313155307290757e+17, 1.31315530739857e+17, 1.313155307507945e+17, 1.313155307611069e+17, 1.313155307712632e+17, 1.313155307817321e+17, 1.313155307918883e+17, 1.313155308025133e+17, 1.313155308128257e+17, 1.313155308237632e+17, 1.313155308339195e+17, 1.313155308440758e+17, 1.313155308543882e+17, 1.313155308648571e+17, 1.313155308751695e+17, 1.313155308868882e+17, 1.313155308976695e+17, 1.313155309078257e+17, 1.313155309181382e+17, 1.313155309287633e+17, 1.313155309395446e+17, 1.31315530949857e+17, 1.313155309600132e+17, 1.313155309703256e+17, 1.313155309812632e+17, 1.313155309915757e+17, 1.313155310028257e+17, 1.31315531012982e+17, 1.313155310239195e+17, 1.31315531034857e+17, 1.313155310451695e+17, 1.313155310557946e+17, 1.313155310664195e+17, 1.313155310770445e+17, 1.313155310876695e+17, 1.313155310981384e+17, 1.313155311082944e+17, 1.31315531118607e+17, 1.31315531129232e+17, 1.313155311397007e+17, 1.313155311506382e+17, 1.313155311611069e+17, 1.31315531171732e+17, 1.313155311826696e+17, 1.31315531193607e+17, 1.313155312040758e+17, 1.313155312143882e+17, 1.31315531224857e+17, 1.313155312350132e+17, 1.313155312451695e+17, 1.313155312553257e+17, 1.313155312659507e+17, 1.313155312764195e+17, 1.313155312870446e+17, 1.313155312975132e+17, 1.313155313076695e+17, 1.313155313179821e+17, 1.313155313282945e+17, 1.31315531339232e+17, 1.313155313500132e+17, 1.313155313601695e+17, 1.31315531370482e+17, 1.313155313807945e+17, 1.313155313912632e+17, 1.313155314028257e+17, 1.313155314131382e+17, 1.313155314232945e+17, 1.313155314337632e+17, 1.313155314445445e+17, 1.31315531454857e+17, 1.313155314651695e+17, 1.313155314756383e+17, 1.313155314864195e+17, 1.313155314965757e+17, 1.313155315068882e+17, 1.313155315173571e+17},
			             {1.313155151125133e+17, 1.313155151226696e+17, 1.31315515132982e+17, 1.313155151434508e+17, 1.313155151550132e+17, 1.313155151653257e+17, 1.31315515175482e+17, 1.313155151857946e+17, 1.313155151959507e+17, 1.313155152065757e+17, 1.313155152175132e+17, 1.31315515227982e+17, 1.313155152382945e+17, 1.313155152487633e+17, 1.313155152593883e+17, 1.313155152700132e+17, 1.313155152807945e+17, 1.313155152911069e+17, 1.313155153022007e+17, 1.313155153126696e+17, 1.313155153232945e+17, 1.313155153334508e+17, 1.313155153439195e+17, 1.313155153542319e+17, 1.31315515364857e+17, 1.313155153751695e+17, 1.313155153856383e+17, 1.313155153957944e+17, 1.31315515406107e+17, 1.313155154173571e+17, 1.313155154281382e+17, 1.313155154390758e+17, 1.313155154501695e+17, 1.31315515460482e+17, 1.31315515471732e+17, 1.313155154825133e+17, 1.313155154926696e+17, 1.313155155032945e+17, 1.313155155134508e+17, 1.313155155240758e+17, 1.31315515534857e+17, 1.313155155451695e+17, 1.313155155559507e+17, 1.313155155665757e+17, 1.313155155765757e+17, 1.313155155875132e+17, 1.313155155976695e+17, 1.313155156078258e+17, 1.313155156184508e+17, 1.313155156293883e+17, 1.313155156397007e+17, 1.313155156501695e+17, 1.313155156607945e+17, 1.313155156714195e+17, 1.313155156818883e+17, 1.313155156928257e+17, 1.31315515702982e+17, 1.313155157131383e+17, 1.31315515723607e+17, 1.313155157340758e+17, 1.313155157442321e+17, 1.313155157543884e+17, 1.313155157651695e+17, 1.313155157757946e+17, 1.31315515786732e+17, 1.313155157968883e+17, 1.313155158072008e+17, 1.313155158173569e+17, 1.313155158275132e+17, 1.313155158376695e+17, 1.313155158479821e+17, 1.31315515857982e+17, 1.313155158681382e+17, 1.313155158789196e+17, 1.313155158890757e+17, 1.313155158995444e+17, 1.313155159103258e+17, 1.313155159211069e+17, 1.313155159312632e+17, 1.313155159414195e+17, 1.31315515952357e+17, 1.313155159625133e+17, 1.31315515972982e+17, 1.31315515982982e+17, 1.313155159931383e+17, 1.313155160039195e+17, 1.31315516014857e+17, 1.313155160251695e+17, 1.31315516035482e+17, 1.31315516046107e+17, 1.313155160565757e+17, 1.313155160668883e+17, 1.313155160776695e+17, 1.313155160881382e+17, 1.313155160984508e+17, 1.313155161086071e+17, 1.31315516119232e+17, 1.31315516129857e+17, 1.313155161411069e+17, 1.313155161522008e+17, 1.313155161625133e+17, 1.313155161728257e+17, 1.313155161831383e+17, 1.313155161937633e+17, 1.313155162039196e+17, 1.313155162143882e+17, 1.313155162247008e+17, 1.313155162356383e+17, 1.313155162462632e+17, 1.31315516256732e+17, 1.313155162668882e+17, 1.313155162772008e+17, 1.313155162875132e+17, 1.313155162978257e+17, 1.313155163081382e+17, 1.313155163182945e+17, 1.313155163284508e+17, 1.31315516339232e+17, 1.313155163501695e+17, 1.313155163603258e+17, 1.313155163706382e+17, 1.313155163811069e+17, 1.313155163912632e+17, 1.313155164014195e+17, 1.313155164115758e+17, 1.313155164215758e+17, 1.313155164326694e+17, 1.313155164428257e+17, 1.313155164531383e+17, 1.313155164639196e+17, 1.313155164745445e+17, 1.313155164847008e+17, 1.313155164953257e+17, 1.313155165062632e+17, 1.313155165164195e+17, 1.313155165270445e+17, 1.313155165375132e+17, 1.313155165478258e+17, 1.313155165581384e+17, 1.313155165684508e+17, 1.313155165787633e+17, 1.31315516589232e+17, 1.313155165993883e+17, 1.313155166097007e+17, 1.313155166200133e+17, 1.31315516630482e+17, 1.313155166409508e+17, 1.313155166514194e+17, 1.313155166615757e+17, 1.313155166718883e+17, 1.313155166831383e+17, 1.31315516693607e+17, 1.313155167045445e+17, 1.313155167150132e+17, 1.313155167253257e+17, 1.313155167362633e+17, 1.313155167462632e+17, 1.313155167564195e+17, 1.313155167675132e+17, 1.313155167784507e+17, 1.31315516788607e+17, 1.313155167989196e+17, 1.31315516809232e+17, 1.313155168195444e+17, 1.313155168297007e+17, 1.313155168403256e+17, 1.31315516850482e+17, 1.313155168612632e+17, 1.313155168714195e+17, 1.313155168820444e+17, 1.313155168922008e+17, 1.313155169037633e+17, 1.313155169143882e+17, 1.313155169245445e+17, 1.313155169351694e+17, 1.31315516945482e+17, 1.313155169568883e+17, 1.313155169672008e+17, 1.313155169776695e+17, 1.313155169887633e+17, 1.31315516999857e+17, 1.313155170101695e+17, 1.31315517020482e+17, 1.313155170307945e+17, 1.313155170411071e+17, 1.313155170514195e+17, 1.313155170618883e+17, 1.313155170720445e+17, 1.313155170822007e+17, 1.313155170931382e+17, 1.313155171037632e+17, 1.313155171139195e+17, 1.313155171242321e+17, 1.313155171343882e+17, 1.313155171447008e+17, 1.313155171551695e+17, 1.31315517166107e+17, 1.313155171765757e+17, 1.313155171868883e+17, 1.313155171970445e+17, 1.313155172170445e+17, 1.313155172278257e+17, 1.313155172382944e+17, 1.313155172484508e+17, 1.313155172589194e+17, 1.313155172693883e+17, 1.313155172795444e+17, 1.313155172900132e+17, 1.313155173006382e+17, 1.313155173109508e+17, 1.313155173214195e+17, 1.313155173315757e+17, 1.313155173418883e+17, 1.31315517352357e+17, 1.313155173626694e+17, 1.31315517372982e+17, 1.313155173832945e+17, 1.31315517393607e+17, 1.313155174039195e+17, 1.313155174142321e+17, 1.313155174243884e+17, 1.313155174347008e+17, 1.31315517444857e+17, 1.313155174551694e+17, 1.313155174653257e+17, 1.313155174757944e+17, 1.313155174865757e+17, 1.313155174978258e+17, 1.313155175082945e+17, 1.313155175193883e+17, 1.31315517529857e+17, 1.31315517540482e+17, 1.313155175507945e+17, 1.31315517562357e+17, 1.313155175725133e+17, 1.313155175837632e+17, 1.313155175940758e+17, 1.313155176042321e+17, 1.313155176143882e+17, 1.313155176243882e+17, 1.313155176345445e+17, 1.313155176453257e+17, 1.31315517656107e+17, 1.313155176665756e+17, 1.313155176768882e+17, 1.313155176872008e+17, 1.313155176973571e+17, 1.31315517707982e+17, 1.313155177184508e+17, 1.313155177290757e+17, 1.313155177395444e+17, 1.31315517749857e+17, 1.313155177600133e+17, 1.313155177704819e+17, 1.313155177807945e+17, 1.313155177912632e+17, 1.313155178017321e+17, 1.313155178122007e+17, 1.31315517822357e+17, 1.313155178325133e+17, 1.31315517842982e+17, 1.313155178534508e+17, 1.313155178639195e+17, 1.313155178747008e+17, 1.313155178850132e+17, 1.313155178959508e+17, 1.31315517906107e+17, 1.313155179165757e+17, 1.313155179273571e+17, 1.313155179375132e+17, 1.313155179482945e+17, 1.31315517958607e+17, 1.313155179687633e+17, 1.313155179793883e+17, 1.313155179895444e+17, 1.31315517999857e+17, 1.31315518009857e+17, 1.313155180200133e+17, 1.313155180307945e+17, 1.313155180411071e+17, 1.313155180514195e+17, 1.313155180617321e+17, 1.313155180718883e+17, 1.313155180822007e+17, 1.31315518092357e+17, 1.313155181028257e+17, 1.31315518112982e+17, 1.313155181232945e+17, 1.313155181340758e+17, 1.313155181442321e+17, 1.313155181543882e+17, 1.313155181645445e+17, 1.313155181753257e+17, 1.31315518185482e+17, 1.313155181957944e+17, 1.313155182065757e+17, 1.313155182172008e+17, 1.313155182273569e+17, 1.31315518237982e+17, 1.31315518247982e+17, 1.313155182584508e+17, 1.313155182695444e+17, 1.313155182801695e+17, 1.313155182904819e+17, 1.313155183012632e+17, 1.313155183115757e+17, 1.31315518322357e+17, 1.313155183325133e+17, 1.313155183428257e+17, 1.313155183531382e+17, 1.313155183634508e+17, 1.313155183747008e+17, 1.31315518386107e+17, 1.31315518396732e+17, 1.313155184075132e+17, 1.31315518417982e+17, 1.313155184284507e+17, 1.31315518438607e+17, 1.313155184492321e+17, 1.313155184595446e+17, 1.31315518469857e+17, 1.313155184801695e+17, 1.313155184907945e+17, 1.313155185014195e+17, 1.313155185122007e+17, 1.313155185226696e+17, 1.313155185326696e+17, 1.313155185439195e+17, 1.313155185545445e+17, 1.313155185645445e+17, 1.31315518575482e+17, 1.313155185856383e+17, 1.313155185959507e+17, 1.31315518606107e+17, 1.313155186173569e+17, 1.313155186276695e+17, 1.313155186378257e+17, 1.31315518648607e+17, 1.313155186595446e+17, 1.313155186701695e+17, 1.313155186806383e+17, 1.313155186909508e+17, 1.313155187011069e+17, 1.313155187115757e+17, 1.31315518721732e+17, 1.313155187318883e+17, 1.31315518742357e+17, 1.313155187525133e+17, 1.313155187628257e+17, 1.313155187739195e+17, 1.313155187840758e+17, 1.313155187945445e+17, 1.313155188047008e+17, 1.313155188150132e+17, 1.313155188253258e+17, 1.31315518836732e+17, 1.313155188476695e+17, 1.313155188578257e+17, 1.31315518867982e+17, 1.313155188782945e+17, 1.313155188884508e+17, 1.313155188987633e+17, 1.313155189090757e+17, 1.313155189195446e+17, 1.313155189303258e+17, 1.31315518940482e+17, 1.313155189506383e+17, 1.313155189607945e+17, 1.313155189714195e+17, 1.313155189815758e+17, 1.313155189918883e+17, 1.31315519002357e+17, 1.313155190126696e+17, 1.313155190232946e+17, 1.31315519033607e+17, 1.313155190439195e+17, 1.313155190542321e+17, 1.31315519064857e+17, 1.313155190750132e+17, 1.313155190850132e+17, 1.313155190953257e+17, 1.313155191059508e+17, 1.31315519116107e+17, 1.313155191264195e+17, 1.313155191365757e+17, 1.31315519146732e+17, 1.313155191570445e+17, 1.313155191681382e+17, 1.313155191784508e+17, 1.313155191887633e+17, 1.313155191987633e+17, 1.313155192089196e+17, 1.313155192195446e+17, 1.31315519229857e+17, 1.31315519240482e+17, 1.313155192506383e+17, 1.313155192612632e+17, 1.313155192714195e+17, 1.31315519281732e+17, 1.313155192920444e+17, 1.313155193026694e+17, 1.313155193126696e+17, 1.31315519323607e+17, 1.313155193340758e+17, 1.313155193445444e+17, 1.313155193550132e+17, 1.31315519365482e+17, 1.313155193757946e+17, 1.31315519386107e+17, 1.313155193964196e+17, 1.31315519406732e+17, 1.313155194168882e+17, 1.313155194273571e+17, 1.313155194376695e+17, 1.313155194484507e+17, 1.313155194590757e+17, 1.31315519469232e+17, 1.313155194800132e+17, 1.313155194901695e+17, 1.31315519500482e+17, 1.313155195106383e+17, 1.313155195211069e+17, 1.31315519531732e+17, 1.313155195418883e+17, 1.31315519552357e+17, 1.313155195625133e+17, 1.313155195726696e+17, 1.313155195832945e+17, 1.313155195940758e+17, 1.31315519605482e+17, 1.313155196157944e+17, 1.31315519626107e+17, 1.313155196372008e+17, 1.313155196476695e+17, 1.31315519657982e+17, 1.313155196681382e+17, 1.31315519678607e+17, 1.313155196889196e+17, 1.313155196989196e+17, 1.313155197093883e+17, 1.313155197203258e+17, 1.31315519730482e+17, 1.313155197409508e+17, 1.313155197512632e+17, 1.31315519761732e+17, 1.313155197720444e+17, 1.313155197825133e+17, 1.313155197926696e+17, 1.313155198032945e+17, 1.313155198140758e+17, 1.313155198242321e+17, 1.313155198345445e+17, 1.313155198450132e+17, 1.31315519855482e+17, 1.31315519866107e+17, 1.31315519876732e+17, 1.313155198878258e+17, 1.313155198984507e+17, 1.313155199089194e+17, 1.313155199195446e+17, 1.313155199306382e+17, 1.313155199420445e+17, 1.313155199522008e+17, 1.31315519962357e+17, 1.313155199726694e+17, 1.313155199828257e+17, 1.31315519992982e+17, 1.313155200037632e+17, 1.313155200150132e+17, 1.313155200251695e+17, 1.313155200353257e+17, 1.313155200456383e+17, 1.313155200562633e+17, 1.313155200664196e+17, 1.313155200772006e+17, 1.31315520087982e+17, 1.31315520098607e+17, 1.31315520109232e+17, 1.313155201193883e+17, 1.313155201297007e+17, 1.31315520140482e+17, 1.313155201506382e+17, 1.313155201607945e+17, 1.313155201714195e+17, 1.313155201822007e+17, 1.313155201925133e+17, 1.313155202026696e+17, 1.313155202134508e+17, 1.313155202236069e+17, 1.313155202337632e+17, 1.313155202439195e+17, 1.313155202550132e+17, 1.313155202653257e+17, 1.313155202754821e+17, 1.313155202868883e+17, 1.313155202972008e+17, 1.313155203073569e+17, 1.313155203178258e+17, 1.313155203282945e+17, 1.31315520339232e+17, 1.313155203495444e+17, 1.31315520359857e+17, 1.313155203704819e+17, 1.313155203811071e+17, 1.313155203914195e+17, 1.313155204014195e+17, 1.313155204115757e+17, 1.313155204225133e+17, 1.313155204326696e+17, 1.313155204437633e+17, 1.313155204540758e+17, 1.313155204643884e+17, 1.313155204750132e+17, 1.313155204850132e+17, 1.313155204953258e+17, 1.313155205057944e+17, 1.313155205162633e+17, 1.313155205264196e+17, 1.313155205365757e+17, 1.313155205468883e+17, 1.313155205570445e+17, 1.313155205676695e+17, 1.313155205789196e+17, 1.313155205900133e+17, 1.31315520600482e+17, 1.313155206112632e+17, 1.313155206215757e+17, 1.313155206318883e+17, 1.313155206422007e+17, 1.313155206526696e+17, 1.31315520663607e+17, 1.313155206743882e+17, 1.313155206847007e+17, 1.313155206951695e+17, 1.313155207057944e+17, 1.313155207165757e+17, 1.313155207270445e+17, 1.31315520737982e+17, 1.31315520748607e+17, 1.313155207587633e+17, 1.313155207689196e+17, 1.313155207793882e+17, 1.313155207900133e+17, 1.313155208007945e+17, 1.313155208112634e+17, 1.31315520821732e+17, 1.313155208326696e+17, 1.31315520842982e+17, 1.31315520852982e+17, 1.313155208634508e+17, 1.313155208740756e+17, 1.313155208842321e+17, 1.313155208943882e+17, 1.313155209047008e+17, 1.313155209150132e+17, 1.313155209253257e+17, 1.31315520936107e+17, 1.31315520946732e+17, 1.313155209575132e+17, 1.313155209675133e+17, 1.313155209781382e+17, 1.31315520988607e+17, 1.313155209997007e+17, 1.313155210107945e+17, 1.313155210211069e+17, 1.313155210311071e+17, 1.313155210412632e+17, 1.313155210514195e+17, 1.31315521061732e+17, 1.31315521072357e+17, 1.313155210826694e+17, 1.31315521092982e+17, 1.313155211037632e+17, 1.313155211140758e+17, 1.313155211248571e+17, 1.31315521136107e+17, 1.31315521146732e+17, 1.313155211568883e+17, 1.313155211672008e+17, 1.313155211773569e+17, 1.313155211878258e+17, 1.313155211982945e+17, 1.313155212087633e+17, 1.313155212200133e+17, 1.31315521230482e+17, 1.313155212407945e+17, 1.313155212511071e+17, 1.313155212622007e+17, 1.313155212725133e+17, 1.313155212839196e+17, 1.313155212943882e+17, 1.31315521304857e+17, 1.313155213153257e+17, 1.31315521325482e+17, 1.313155213357944e+17, 1.31315521346107e+17, 1.31315521356732e+17, 1.313155213678258e+17, 1.313155213781382e+17, 1.313155213884508e+17, 1.31315521398607e+17, 1.313155214087633e+17, 1.313155214287633e+17, 1.313155214393883e+17, 1.313155214500132e+17, 1.313155214609508e+17, 1.313155214712632e+17, 1.313155214815757e+17, 1.313155214918883e+17, 1.313155215022007e+17, 1.31315521512357e+17, 1.313155215226696e+17, 1.31315521533607e+17, 1.313155215439196e+17, 1.313155215547007e+17, 1.31315521564857e+17, 1.313155215764195e+17, 1.31315521586732e+17, 1.313155215976695e+17, 1.31315521607982e+17, 1.313155216182945e+17, 1.313155216287631e+17, 1.313155216389194e+17, 1.31315521649232e+17, 1.313155216595444e+17, 1.313155216700132e+17, 1.313155216807945e+17, 1.313155216912632e+17, 1.313155217012634e+17, 1.313155217115758e+17, 1.313155217218883e+17, 1.313155217325133e+17, 1.313155217434508e+17, 1.31315521753607e+17, 1.31315521764857e+17, 1.313155217750132e+17, 1.313155217851695e+17, 1.313155217953258e+17, 1.31315521805482e+17, 1.313155218159507e+17, 1.31315521826107e+17, 1.313155218362633e+17, 1.313155218465757e+17, 1.313155218578257e+17, 1.313155218682945e+17, 1.313155218789196e+17, 1.313155218897007e+17, 1.31315521899857e+17, 1.313155219101696e+17, 1.313155219212632e+17, 1.313155219315757e+17, 1.313155219418883e+17, 1.31315521952357e+17, 1.313155219626694e+17, 1.313155219737632e+17, 1.313155219839195e+17, 1.313155219939195e+17, 1.313155220040758e+17, 1.313155220143882e+17, 1.313155220250134e+17, 1.313155220351695e+17, 1.313155220453257e+17, 1.313155220556383e+17, 1.31315522066107e+17, 1.313155220764195e+17, 1.313155220867319e+17, 1.313155220968882e+17, 1.313155221075132e+17, 1.313155221182944e+17, 1.313155221293883e+17, 1.313155221401695e+17, 1.313155221509508e+17, 1.313155221611071e+17, 1.31315522171732e+17, 1.313155221828257e+17, 1.31315522192982e+17, 1.313155222039195e+17, 1.313155222140758e+17, 1.313155222245445e+17, 1.313155222353258e+17, 1.313155222464195e+17, 1.31315522256732e+17, 1.313155222672006e+17, 1.313155222773569e+17, 1.313155222875132e+17, 1.313155222989196e+17, 1.313155223097007e+17, 1.31315522319857e+17, 1.313155223303256e+17, 1.31315522340482e+17, 1.313155223511069e+17, 1.313155223612632e+17, 1.313155223714195e+17, 1.313155223820444e+17, 1.313155223920445e+17, 1.31315522402982e+17, 1.31315522413607e+17, 1.313155224237633e+17, 1.313155224342319e+17, 1.313155224442321e+17, 1.31315522454857e+17, 1.313155224650132e+17, 1.313155224751695e+17, 1.31315522485482e+17, 1.313155224957946e+17, 1.31315522506107e+17, 1.313155225162633e+17, 1.313155225264196e+17, 1.31315522536732e+17, 1.313155225470445e+17, 1.313155225578258e+17, 1.313155225682945e+17, 1.313155225784508e+17, 1.313155225887633e+17, 1.313155225993883e+17, 1.313155226104819e+17, 1.313155226214194e+17, 1.31315522631732e+17, 1.313155226420444e+17, 1.31315522652357e+17, 1.313155226628257e+17, 1.313155226742319e+17, 1.313155226843882e+17, 1.313155226945445e+17, 1.313155227047007e+17, 1.31315522714857e+17, 1.313155227253257e+17, 1.313155227359507e+17, 1.313155227462633e+17, 1.313155227564196e+17, 1.313155227668883e+17, 1.313155227773571e+17, 1.313155227876695e+17, 1.313155227984508e+17, 1.31315522808607e+17, 1.313155228193882e+17, 1.313155228295444e+17, 1.31315522839857e+17, 1.313155228503258e+17, 1.313155228612632e+17, 1.313155228726696e+17, 1.313155228831382e+17, 1.313155228934508e+17, 1.313155229045445e+17, 1.313155229151695e+17, 1.313155229262633e+17, 1.313155229365757e+17, 1.31315522947982e+17, 1.313155229584508e+17, 1.313155229690758e+17, 1.313155229804819e+17, 1.313155229911071e+17, 1.313155230022007e+17, 1.31315523012357e+17, 1.313155230228257e+17, 1.31315523032982e+17, 1.313155230431383e+17, 1.313155230534508e+17, 1.313155230642319e+17, 1.313155230743882e+17, 1.313155230847008e+17, 1.313155230953257e+17, 1.31315523105482e+17, 1.313155231156383e+17, 1.313155231270445e+17, 1.313155231379821e+17, 1.313155231484508e+17, 1.313155231592321e+17, 1.31315523169857e+17, 1.313155231801695e+17, 1.313155231906382e+17, 1.313155232011071e+17, 1.313155232114195e+17, 1.313155232214195e+17, 1.313155232318883e+17, 1.313155232418883e+17, 1.313155232525133e+17, 1.313155232634508e+17, 1.313155232739195e+17, 1.313155232842319e+17, 1.313155232945445e+17, 1.31315523304857e+17, 1.313155233150132e+17, 1.313155233251695e+17, 1.313155233353257e+17, 1.31315523345482e+17, 1.313155233556383e+17, 1.31315523366107e+17, 1.313155233764195e+17, 1.313155233865757e+17, 1.313155233973571e+17, 1.313155234078258e+17, 1.313155234179821e+17, 1.31315523428607e+17, 1.313155234390757e+17, 1.31315523449232e+17, 1.31315523459232e+17, 1.31315523469857e+17, 1.313155234800133e+17, 1.313155234911069e+17, 1.313155235014195e+17, 1.313155235126694e+17, 1.313155235236069e+17, 1.313155235343882e+17, 1.31315523544857e+17, 1.313155235556383e+17, 1.313155235657946e+17, 1.313155235765757e+17, 1.313155235870445e+17, 1.313155235975132e+17, 1.313155236081382e+17, 1.31315523618607e+17, 1.313155236289196e+17, 1.31315523639232e+17, 1.313155236593883e+17, 1.313155236695446e+17, 1.313155236797007e+17, 1.313155236900132e+17, 1.313155237003256e+17, 1.313155237106382e+17, 1.313155237209508e+17, 1.313155237309508e+17, 1.313155237414195e+17, 1.313155237515758e+17, 1.313155237618883e+17, 1.313155237720444e+17, 1.313155237825133e+17, 1.313155237928257e+17, 1.313155238037633e+17, 1.313155238142321e+17, 1.313155238243882e+17, 1.313155238345444e+17, 1.313155238447008e+17, 1.313155238548571e+17, 1.313155238653257e+17, 1.313155238765757e+17, 1.31315523886732e+17, 1.313155238976695e+17, 1.313155239078258e+17, 1.313155239187633e+17, 1.313155239297007e+17, 1.313155239400133e+17, 1.313155239514195e+17, 1.313155239615757e+17, 1.313155239725133e+17, 1.31315523982982e+17, 1.313155239934508e+17, 1.313155240037633e+17, 1.313155240142321e+17, 1.31315524025482e+17, 1.313155240359507e+17, 1.313155240462633e+17, 1.313155240570445e+17, 1.313155240675132e+17, 1.31315524078607e+17, 1.31315524089232e+17, 1.31315524099232e+17, 1.313155241095444e+17, 1.31315524119857e+17, 1.313155241301695e+17, 1.313155241406382e+17, 1.313155241507945e+17, 1.313155241609508e+17, 1.313155241714195e+17, 1.313155241815758e+17, 1.313155241926696e+17, 1.313155242032945e+17, 1.313155242134508e+17, 1.313155242242321e+17, 1.313155242345445e+17, 1.313155242450132e+17, 1.313155242551695e+17, 1.313155242657944e+17, 1.31315524276732e+17, 1.313155242870445e+17, 1.313155242978258e+17, 1.313155243090757e+17, 1.313155243193883e+17, 1.313155243301695e+17, 1.313155243406382e+17, 1.313155243514195e+17, 1.313155243615758e+17, 1.313155243715757e+17, 1.313155243818883e+17, 1.313155243922007e+17, 1.313155244025133e+17, 1.313155244139195e+17, 1.313155244240758e+17, 1.31315524434857e+17, 1.313155244451695e+17, 1.313155244553257e+17, 1.313155244656383e+17, 1.31315524476107e+17, 1.313155244862633e+17, 1.313155244973569e+17, 1.313155245082944e+17, 1.313155245184508e+17, 1.313155245286071e+17, 1.313155245395444e+17, 1.313155245501695e+17, 1.313155245609508e+17, 1.313155245718883e+17, 1.31315524582357e+17, 1.313155245928257e+17, 1.313155246032945e+17, 1.313155246134508e+17, 1.31315524623607e+17, 1.313155246340756e+17, 1.313155246442321e+17, 1.313155246543884e+17, 1.313155246647008e+17, 1.313155246750132e+17, 1.313155246857944e+17, 1.31315524696107e+17, 1.31315524706732e+17, 1.313155247168883e+17, 1.313155247281382e+17, 1.31315524738607e+17, 1.313155247489194e+17, 1.313155247603258e+17, 1.313155247711071e+17, 1.31315524781732e+17, 1.313155247922008e+17, 1.313155248028257e+17, 1.31315524813607e+17, 1.313155248239195e+17, 1.313155248340758e+17, 1.313155248445445e+17, 1.31315524855482e+17, 1.313155248657946e+17, 1.313155248762633e+17, 1.313155248870445e+17, 1.313155248973571e+17, 1.313155249075132e+17, 1.313155249178257e+17, 1.313155249282945e+17, 1.313155249392321e+17, 1.313155249493883e+17, 1.31315524959857e+17, 1.313155249700132e+17, 1.313155249803258e+17, 1.313155249912632e+17, 1.313155250022007e+17, 1.313155250126696e+17, 1.313155250232945e+17, 1.31315525033607e+17, 1.313155250437633e+17, 1.313155250543882e+17, 1.313155250645445e+17, 1.31315525074857e+17, 1.31315525085482e+17, 1.313155250962632e+17, 1.313155251064195e+17, 1.313155251165757e+17, 1.313155251265757e+17, 1.313155251370445e+17, 1.313155251476695e+17, 1.313155251586071e+17, 1.313155251690757e+17, 1.31315525179232e+17, 1.313155251893882e+17, 1.313155251997007e+17, 1.313155252100132e+17, 1.313155252201695e+17, 1.313155252311069e+17, 1.313155252415757e+17, 1.313155252520445e+17, 1.31315525262357e+17, 1.313155252734508e+17, 1.313155252843884e+17, 1.313155252947008e+17, 1.31315525304857e+17, 1.313155253153258e+17, 1.313155253259507e+17, 1.31315525336732e+17, 1.313155253470445e+17, 1.313155253572008e+17, 1.313155253676695e+17, 1.313155253784508e+17, 1.31315525388607e+17, 1.313155254001695e+17, 1.313155254106383e+17, 1.313155254206382e+17, 1.313155254311069e+17, 1.313155254414194e+17, 1.313155254518883e+17, 1.31315525462357e+17, 1.313155254726696e+17, 1.313155254831383e+17, 1.313155254934508e+17, 1.313155255037633e+17, 1.313155255142319e+17, 1.313155255243882e+17, 1.313155255345445e+17, 1.31315525545482e+17, 1.313155255559507e+17, 1.313155255664195e+17, 1.31315525576732e+17, 1.313155255868883e+17, 1.313155255970445e+17, 1.313155256073569e+17, 1.313155256176695e+17, 1.313155256278258e+17, 1.313155256382944e+17, 1.313155256484507e+17, 1.31315525658607e+17, 1.313155256693883e+17, 1.31315525679857e+17, 1.313155256900133e+17, 1.313155257006383e+17, 1.313155257109508e+17, 1.313155257212632e+17, 1.313155257314195e+17, 1.313155257417321e+17, 1.31315525752357e+17, 1.313155257628257e+17, 1.313155257734508e+17, 1.313155257842321e+17, 1.313155257951695e+17, 1.313155258053257e+17, 1.31315525815482e+17, 1.313155258257946e+17, 1.313155258370445e+17, 1.313155258475132e+17, 1.313155258579821e+17, 1.313155258682945e+17, 1.31315525879232e+17, 1.31315525889857e+17, 1.313155259003258e+17, 1.313155259103258e+17, 1.313155259206382e+17, 1.313155259311069e+17, 1.313155259412632e+17, 1.31315525952357e+17, 1.313155259632945e+17, 1.31315525973607e+17, 1.313155259837633e+17, 1.313155259942319e+17, 1.313155260043882e+17, 1.313155260145445e+17, 1.313155260250132e+17, 1.313155260353257e+17, 1.313155260457944e+17, 1.31315526056107e+17, 1.313155260665757e+17, 1.313155260773571e+17, 1.313155260875133e+17, 1.313155260982945e+17, 1.313155261095444e+17, 1.31315526119857e+17, 1.31315526130482e+17, 1.313155261407945e+17, 1.313155261509507e+17, 1.313155261611069e+17, 1.313155261714195e+17, 1.313155261825133e+17, 1.31315526192982e+17, 1.313155262031383e+17, 1.313155262134508e+17, 1.313155262240758e+17, 1.313155262359507e+17, 1.31315526246107e+17, 1.313155262564195e+17, 1.31315526266732e+17, 1.31315526277982e+17, 1.313155262882944e+17, 1.31315526298607e+17, 1.31315526309232e+17, 1.313155263193883e+17, 1.313155263297007e+17, 1.313155263400132e+17, 1.313155263506382e+17, 1.313155263611069e+17, 1.313155263712632e+17, 1.313155263815757e+17, 1.313155263926696e+17, 1.31315526402982e+17, 1.313155264132945e+17, 1.31315526423607e+17, 1.313155264337633e+17, 1.313155264445445e+17, 1.31315526454857e+17, 1.313155264657946e+17, 1.31315526476107e+17, 1.313155264864195e+17, 1.313155264970445e+17, 1.313155265073571e+17, 1.313155265181382e+17, 1.313155265287633e+17, 1.313155265395444e+17, 1.313155265509508e+17, 1.313155265611069e+17, 1.313155265715758e+17, 1.313155265822007e+17, 1.313155265925133e+17, 1.313155266037633e+17, 1.313155266140758e+17, 1.313155266243882e+17, 1.313155266347008e+17, 1.31315526644857e+17, 1.313155266553257e+17, 1.313155266659507e+17, 1.31315526676107e+17, 1.313155266864196e+17, 1.313155266973571e+17, 1.313155267078258e+17, 1.313155267184507e+17, 1.313155267290757e+17, 1.31315526740482e+17, 1.313155267507945e+17, 1.313155267618883e+17, 1.313155267720445e+17, 1.31315526782357e+17, 1.313155267925133e+17, 1.313155268032945e+17, 1.31315526813607e+17, 1.313155268237633e+17, 1.313155268339195e+17, 1.313155268442319e+17, 1.31315526855482e+17, 1.313155268672008e+17, 1.31315526877982e+17, 1.31315526888607e+17, 1.31315526899232e+17, 1.313155269093883e+17, 1.31315526919857e+17, 1.313155269301696e+17, 1.31315526940482e+17, 1.313155269507945e+17, 1.313155269609508e+17, 1.313155269712632e+17, 1.31315526982982e+17, 1.313155269936069e+17, 1.313155270045445e+17, 1.31315527014857e+17, 1.313155270257944e+17, 1.313155270359507e+17, 1.313155270462633e+17, 1.313155270565757e+17, 1.313155270673571e+17, 1.313155270778258e+17, 1.313155270882944e+17, 1.31315527098607e+17, 1.313155271087633e+17, 1.31315527119232e+17, 1.313155271295444e+17, 1.313155271400132e+17, 1.313155271506383e+17, 1.313155271614195e+17, 1.313155271715757e+17, 1.313155271822008e+17, 1.31315527193607e+17, 1.313155272042321e+17, 1.313155272147007e+17, 1.313155272250132e+17, 1.313155272353257e+17, 1.31315527245482e+17, 1.313155272557944e+17, 1.31315527266107e+17, 1.313155272764196e+17, 1.313155272873571e+17, 1.313155272976695e+17, 1.313155273082944e+17, 1.313155273184507e+17, 1.313155273290757e+17, 1.313155273395446e+17, 1.313155273501695e+17, 1.313155273603258e+17, 1.313155273706383e+17, 1.313155273809508e+17, 1.313155273911071e+17, 1.31315527401732e+17, 1.31315527412357e+17, 1.313155274225133e+17, 1.313155274331383e+17, 1.313155274431382e+17, 1.313155274540758e+17, 1.313155274642321e+17, 1.313155274745445e+17, 1.313155274845445e+17, 1.313155274959507e+17, 1.31315527506107e+17, 1.313155275162633e+17, 1.313155275265757e+17, 1.313155275367319e+17, 1.313155275472008e+17, 1.313155275575132e+17, 1.313155275679821e+17, 1.313155275782945e+17, 1.313155275897007e+17, 1.313155276003258e+17, 1.313155276114195e+17, 1.31315527622357e+17, 1.313155276323571e+17, 1.31315527643607e+17, 1.313155276539195e+17, 1.313155276642319e+17, 1.313155276745445e+17, 1.313155276851695e+17, 1.31315527696107e+17, 1.313155277062632e+17, 1.313155277165757e+17, 1.31315527726732e+17, 1.313155277368883e+17, 1.313155277476695e+17, 1.31315527758607e+17, 1.313155277690757e+17, 1.313155277800133e+17, 1.313155277903258e+17, 1.31315527801732e+17, 1.313155278126696e+17, 1.313155278237633e+17, 1.313155278340758e+17, 1.313155278450132e+17, 1.31315527856107e+17, 1.31315527866732e+17, 1.313155278778258e+17, 1.313155278884507e+17, 1.313155278989196e+17, 1.313155279093883e+17, 1.313155279195444e+17, 1.313155279301695e+17, 1.313155279403258e+17, 1.313155279509508e+17, 1.313155279609508e+17, 1.313155279718883e+17, 1.313155279820444e+17, 1.313155279922007e+17, 1.31315528002357e+17, 1.313155280125133e+17, 1.313155280237633e+17, 1.313155280339196e+17, 1.313155280440758e+17, 1.31315528054857e+17, 1.313155280654821e+17, 1.313155280759507e+17, 1.313155280862633e+17, 1.313155280972008e+17, 1.313155281075132e+17, 1.313155281178258e+17, 1.313155281279821e+17, 1.313155281382945e+17, 1.313155281495444e+17, 1.313155281600132e+17, 1.313155281703258e+17, 1.313155281807945e+17, 1.313155281911069e+17, 1.313155282012632e+17, 1.313155282128257e+17, 1.313155282242319e+17, 1.313155282345445e+17, 1.313155282456383e+17, 1.313155282562633e+17, 1.313155282664195e+17, 1.313155282765757e+17, 1.31315528286732e+17, 1.313155282975133e+17, 1.313155283082944e+17, 1.31315528318607e+17, 1.313155283287633e+17, 1.313155283389196e+17, 1.313155283495444e+17, 1.313155283607945e+17, 1.313155283709508e+17, 1.313155283814195e+17, 1.313155283931383e+17, 1.313155284034508e+17, 1.31315528413607e+17, 1.313155284239195e+17, 1.313155284343882e+17, 1.313155284445445e+17, 1.313155284553257e+17, 1.313155284662632e+17, 1.313155284764195e+17, 1.313155284868882e+17, 1.313155284972006e+17, 1.313155285075132e+17, 1.313155285182945e+17, 1.313155285290757e+17, 1.313155285395444e+17, 1.31315528549857e+17, 1.31315528559857e+17, 1.313155285701695e+17, 1.313155285803258e+17, 1.313155285907945e+17, 1.313155286020444e+17, 1.31315528612357e+17, 1.313155286232945e+17, 1.313155286342321e+17, 1.31315528645482e+17, 1.313155286557944e+17, 1.313155286657944e+17, 1.313155286765757e+17, 1.313155286868883e+17, 1.313155286970445e+17, 1.31315528707982e+17, 1.313155287193883e+17, 1.313155287301695e+17, 1.313155287407944e+17, 1.313155287512632e+17, 1.313155287618883e+17, 1.313155287720445e+17, 1.313155287825133e+17, 1.313155287932945e+17, 1.31315528803607e+17, 1.313155288137632e+17, 1.313155288247007e+17, 1.313155288357946e+17, 1.313155288462633e+17, 1.313155288570445e+17, 1.313155288675133e+17, 1.313155288784508e+17, 1.313155288889196e+17, 1.31315528899857e+17, 1.313155289115757e+17, 1.31315528921732e+17, 1.313155289318883e+17, 1.313155289431382e+17, 1.313155289534508e+17, 1.313155289637632e+17, 1.313155289740756e+17, 1.313155289842321e+17, 1.313155289945445e+17, 1.31315529004857e+17, 1.313155290153257e+17, 1.313155290253258e+17, 1.31315529035482e+17, 1.313155290457944e+17, 1.313155290572008e+17, 1.313155290676695e+17, 1.313155290778258e+17, 1.313155290879821e+17, 1.313155290982945e+17, 1.313155291084507e+17, 1.313155291193883e+17, 1.313155291295444e+17, 1.31315529139857e+17, 1.31315529150482e+17, 1.313155291612632e+17, 1.313155291715757e+17, 1.31315529181732e+17, 1.313155291922007e+17, 1.313155292028257e+17, 1.313155292142321e+17, 1.313155292251695e+17, 1.313155292362633e+17, 1.313155292464196e+17, 1.313155292565757e+17, 1.313155292670445e+17, 1.313155292773571e+17, 1.313155292875132e+17, 1.31315529297982e+17, 1.313155293079821e+17, 1.313155293182945e+17, 1.313155293290757e+17, 1.313155293401695e+17, 1.313155293511069e+17, 1.313155293612632e+17, 1.313155293714194e+17, 1.313155293818883e+17, 1.313155293922008e+17, 1.31315529402357e+17, 1.313155294125133e+17, 1.313155294226696e+17, 1.313155294331383e+17, 1.313155294434508e+17, 1.313155294543882e+17, 1.313155294651695e+17, 1.313155294765757e+17, 1.31315529487982e+17, 1.313155294981382e+17, 1.313155295084507e+17, 1.313155295187633e+17, 1.313155295287631e+17, 1.313155295393883e+17, 1.313155295495446e+17, 1.31315529559857e+17, 1.313155295700132e+17, 1.313155295801695e+17, 1.313155295907945e+17, 1.313155296012634e+17, 1.313155296115758e+17, 1.313155296225133e+17, 1.31315529632982e+17, 1.313155296434508e+17, 1.313155296540758e+17, 1.313155296651695e+17, 1.313155296751695e+17, 1.313155296853257e+17, 1.313155296956383e+17, 1.313155297056383e+17, 1.313155297159507e+17, 1.313155297265757e+17, 1.31315529736732e+17, 1.313155297482945e+17, 1.313155297593883e+17, 1.31315529769857e+17, 1.313155297803258e+17, 1.313155297911069e+17, 1.313155298012632e+17, 1.313155298118883e+17, 1.313155298220444e+17, 1.313155298326696e+17, 1.313155298437633e+17, 1.313155298539195e+17, 1.313155298642321e+17, 1.313155298743882e+17, 1.313155298847007e+17, 1.313155298953257e+17, 1.313155299057946e+17, 1.313155299159508e+17, 1.31315529926107e+17, 1.313155299362633e+17, 1.313155299464196e+17, 1.313155299565757e+17, 1.31315529966732e+17, 1.313155299775132e+17, 1.313155299878257e+17, 1.313155299981382e+17, 1.313155300090757e+17, 1.31315530019857e+17, 1.313155300301695e+17, 1.313155300403258e+17, 1.313155300507945e+17, 1.313155300614195e+17, 1.313155300722008e+17, 1.313155300823571e+17, 1.313155300928257e+17, 1.31315530102982e+17, 1.313155301131382e+17, 1.313155301232945e+17, 1.313155301340758e+17, 1.313155301457944e+17, 1.313155301564195e+17, 1.31315530166732e+17, 1.313155301768882e+17, 1.313155301872008e+17, 1.313155301976695e+17, 1.313155302078257e+17, 1.313155302182944e+17, 1.313155302284508e+17, 1.313155302397009e+17, 1.313155302500133e+17, 1.313155302603258e+17, 1.313155302704819e+17, 1.313155302812632e+17, 1.313155302920445e+17, 1.31315530302357e+17, 1.313155303126696e+17, 1.31315530322982e+17, 1.313155303331382e+17, 1.313155303437632e+17, 1.313155303539195e+17, 1.313155303640756e+17, 1.313155303743882e+17, 1.313155303845445e+17, 1.313155303947008e+17, 1.313155304056383e+17, 1.313155304159507e+17, 1.313155304265757e+17, 1.313155304368882e+17, 1.313155304472008e+17, 1.313155304575132e+17, 1.313155304687633e+17, 1.313155304789194e+17, 1.31315530489232e+17, 1.313155304997007e+17, 1.313155305104819e+17, 1.31315530520482e+17, 1.313155305306382e+17, 1.313155305407945e+17, 1.313155305514195e+17, 1.313155305617321e+17, 1.313155305720445e+17, 1.313155305822007e+17, 1.31315530592357e+17, 1.313155306025133e+17, 1.313155306128257e+17, 1.31315530622982e+17, 1.313155306331382e+17, 1.313155306440758e+17, 1.313155306543882e+17, 1.313155306659507e+17, 1.313155306765757e+17, 1.31315530686732e+17, 1.313155306972008e+17, 1.313155307075133e+17, 1.313155307181382e+17, 1.313155307290757e+17, 1.31315530739857e+17, 1.313155307507945e+17, 1.313155307611069e+17, 1.313155307712632e+17, 1.313155307817321e+17, 1.313155307918883e+17, 1.313155308025133e+17, 1.313155308128257e+17, 1.313155308237632e+17, 1.313155308339195e+17, 1.313155308440758e+17, 1.313155308543882e+17, 1.313155308648571e+17, 1.313155308751695e+17, 1.313155308868882e+17, 1.313155308976695e+17, 1.313155309078257e+17, 1.313155309181382e+17, 1.313155309287633e+17, 1.313155309395446e+17, 1.31315530949857e+17, 1.313155309600132e+17, 1.313155309703256e+17, 1.313155309812632e+17, 1.313155309915757e+17, 1.313155310028257e+17, 1.31315531012982e+17, 1.313155310239195e+17, 1.31315531034857e+17, 1.313155310451695e+17, 1.313155310557946e+17, 1.313155310664195e+17, 1.313155310770445e+17, 1.313155310876695e+17, 1.313155310981384e+17, 1.313155311082944e+17, 1.31315531118607e+17, 1.31315531129232e+17, 1.313155311397007e+17, 1.313155311506382e+17, 1.313155311611069e+17, 1.31315531171732e+17, 1.313155311826696e+17, 1.31315531193607e+17, 1.313155312040758e+17, 1.313155312143882e+17, 1.31315531224857e+17, 1.313155312350132e+17, 1.313155312451695e+17, 1.313155312553257e+17, 1.313155312659507e+17, 1.313155312764195e+17, 1.313155312870446e+17, 1.313155312975132e+17, 1.313155313076695e+17, 1.313155313179821e+17, 1.313155313282945e+17, 1.31315531339232e+17, 1.313155313500132e+17, 1.313155313601695e+17, 1.31315531370482e+17, 1.313155313807945e+17, 1.313155313912632e+17, 1.313155314028257e+17, 1.313155314131382e+17, 1.313155314232945e+17, 1.313155314337632e+17, 1.313155314445445e+17, 1.31315531454857e+17, 1.313155314651695e+17, 1.313155314756383e+17, 1.313155314864195e+17, 1.313155314965757e+17, 1.313155315068882e+17, 1.313155315173571e+17};
			mask_depths = {{15.0, 15.0, 66.8, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 66.8}, {15.0, 15.0, 60.3, 60.3, 66.8, 72.9}}, {{66.8, 66.8, 93.6, 93.6}, {66.8, 93.5}, {66.8, 93.5}, {66.8, 93.3}, {66.8, 93.4}, {66.8, 93.5}, {66.8, 93.7}, {66.8, 93.4}, {66.8, 93.4}, {66.8, 93.4}, {66.8, 93.5}, {66.8, 93.5}, {66.8, 93.4}, {66.8, 93.5}, {66.8, 93.5}, {66.8, 93.4}, {66.8, 93.2}, {66.8, 93.1}, {66.8, 92.9}, {66.8, 92.9}, {66.8, 93.1}, {66.8, 93.3}, {66.8, 93.0}, {66.8, 92.7}, {66.8, 93.2}, {66.8, 93.2}, {66.8, 92.9}, {66.8, 93.1}, {66.8, 93.3}, {66.8, 93.3}, {66.8, 93.5}, {66.8, 93.4}, {66.8, 93.4}, {66.8, 93.4}, {66.8, 93.5}, {66.8, 93.5}, {66.8, 93.7}, {66.8, 93.7}, {66.8, 93.6}, {66.8, 93.6}, {66.8, 93.6}, {66.8, 93.5}, {66.8, 93.4}, {66.8, 93.5}, {66.8, 93.5}, {66.8, 93.4}, {66.8, 93.7}, {66.8, 93.9}, {66.8, 93.9}, {66.8, 93.8}, {66.8, 93.5}, {66.8, 93.6}, {66.8, 93.5}, {66.8, 93.5}, {66.8, 93.6}, {66.8, 93.6}, {66.8, 93.8}, {66.8, 93.9}, {66.8, 94.0}, {66.8, 94.0}, {66.8, 93.9}, {66.8, 93.9}, {66.8, 94.0}, {66.8, 94.1}, {66.8, 94.3}, {66.8, 94.3}, {66.8, 94.2}, {66.8, 94.5}, {66.8, 94.7}, {66.8, 94.5}, {66.8, 94.6}, {66.8, 94.3}, {66.8, 94.5}, {66.8, 94.7}, {66.8, 94.6}, {66.8, 94.8}, {66.8, 94.7}, {66.8, 94.3}, {66.8, 94.8}, {66.8, 94.8}, {66.8, 94.7}, {66.8, 94.6}, {66.8, 94.7}, {66.8, 94.7}, {66.8, 94.6}, {66.8, 94.6}, {66.8, 94.5}, {66.8, 94.4}, {66.8, 94.4}, {66.8, 94.2}, {66.8, 94.3}, {66.8, 94.2}, {66.8, 94.3}, {66.8, 94.4}, {66.8, 94.3}, {66.8, 94.3}, {66.8, 94.3}, {66.8, 94.4}, {66.8, 94.2}, {66.8, 94.2}, {66.8, 94.4}, {66.8, 94.3}, {66.8, 94.4}, {66.8, 94.3}, {66.8, 94.2}, {66.8, 94.4}, {66.8, 94.6}, {66.8, 94.5}, {66.8, 94.6}, {66.8, 94.6}, {66.8, 94.7}, {66.8, 94.6}, {66.8, 94.4}, {66.8, 94.4}, {66.8, 94.5}, {66.8, 94.5}, {66.8, 94.8}, {66.8, 94.9}, {66.8, 94.9}, {66.8, 95.2}, {66.8, 95.0}, {66.8, 95.0}, {66.8, 95.0}, {66.8, 95.2}, {66.8, 95.4}, {66.8, 95.4}, {66.8, 95.4}, {66.8, 95.4}, {66.8, 95.3}, {66.8, 95.3}, {66.8, 95.1}, {66.8, 95.1}, {66.8, 95.3}, {66.8, 95.5}, {66.8, 95.6}, {66.8, 95.6}, {66.8, 95.6}, {66.8, 95.5}, {66.8, 95.5}, {66.8, 95.6}, {66.8, 95.7}, {66.8, 95.6}, {66.8, 95.6}, {66.8, 95.8}, {66.8, 96.1}, {66.8, 96.2}, {66.8, 96.1}, {66.8, 96.4}, {66.8, 96.5}, {66.8, 96.5}, {66.8, 96.3}, {66.8, 96.2}, {66.8, 96.3}, {66.8, 96.3}, {66.8, 96.3}, {66.8, 96.4}, {66.8, 96.3}, {66.8, 96.6}, {66.8, 96.7}, {66.8, 96.7}, {66.8, 96.6}, {66.8, 96.4}, {66.8, 96.2}, {66.8, 96.1}, {66.8, 96.3}, {66.8, 96.3}, {66.8, 96.3}, {66.8, 96.4}, {66.8, 96.3}, {66.8, 96.3}, {66.8, 96.1}, {66.8, 96.0}, {66.8, 96.0}, {66.8, 96.0}, {66.8, 95.8}, {66.8, 95.8}, {66.8, 96.1}, {66.8, 96.1}, {66.8, 96.1}, {66.8, 96.2}, {66.8, 96.2}, {66.8, 96.1}, {66.8, 96.0}, {66.8, 96.2}, {66.8, 96.2}, {66.8, 96.2}, {66.8, 96.3}, {66.8, 96.5}, {66.8, 96.5}, {66.8, 96.5}, {66.8, 96.4}, {66.8, 96.3}, {66.8, 96.3}, {66.8, 96.5}, {66.8, 96.5}, {66.8, 96.8}, {66.8, 96.9}, {66.8, 97.1}, {66.8, 97.1}, {66.8, 96.7}, {66.8, 96.6}, {66.8, 97.0}, {66.8, 96.8}, {66.8, 96.9}, {66.8, 97.1}, {66.8, 97.1}, {66.8, 97.2}, {66.8, 97.1}, {66.8, 97.1}, {66.8, 97.1}, {66.8, 97.3}, {66.8, 97.4}, {66.8, 97.5}, {66.8, 97.4}, {66.8, 97.5}, {66.8, 97.4}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.4}, {66.8, 97.3}, {66.8, 97.4}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.7}, {66.8, 97.6}, {66.8, 97.4}, {66.8, 97.3}, {66.8, 97.4}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.4}, {66.8, 97.6}, {66.8, 97.5}, {66.8, 97.4}, {66.8, 97.4}, {66.8, 97.2}, {66.8, 97.0}, {66.8, 97.0}, {66.8, 96.9}, {66.8, 96.8}, {66.8, 97.0}, {66.8, 97.3}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.2}, {66.8, 96.9}, {66.8, 97.6}, {66.8, 97.7}, {66.8, 97.7}, {66.8, 97.8}, {66.8, 97.8}, {66.8, 97.9}, {66.8, 97.8}, {66.8, 97.7}, {66.8, 97.7}, {66.8, 97.7}, {66.8, 97.6}, {66.8, 97.4}, {66.8, 97.4}, {66.8, 97.8}, {66.8, 97.8}, {66.8, 97.7}, {66.8, 97.8}, {66.8, 97.7}, {66.8, 97.8}, {66.8, 97.8}, {66.8, 97.6}, {66.8, 97.6}, {66.8, 97.4}, {66.8, 96.9}, {66.8, 97.4}, {66.8, 97.4}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.6}, {66.8, 97.7}, {66.8, 97.7}, {66.8, 97.8}, {66.8, 97.9}, {66.8, 97.9}, {66.8, 97.8}, {66.8, 97.4}, {66.8, 97.3}, {66.8, 97.3}, {66.8, 97.5}, {66.8, 97.8}, {66.8, 97.9}, {66.8, 98.1}, {66.8, 98.2}, {66.8, 98.3}, {66.8, 98.3}, {66.8, 98.2}, {66.8, 98.2}, {66.8, 98.0}, {66.8, 97.7}, {66.8, 97.7}, {66.8, 97.7}, {66.8, 97.8}, {66.8, 97.7}, {66.8, 97.6}, {66.8, 97.3}, {66.8, 97.4}, {66.8, 97.4}, {66.8, 97.3}, {66.8, 97.4}, {66.8, 97.3}, {66.8, 97.2}, {66.8, 97.5}, {66.8, 97.5}, {66.8, 97.4}, {66.8, 97.2}, {66.8, 97.3}, {66.8, 97.2}, {66.8, 97.1}, {66.8, 97.1}, {66.8, 97.2}, {66.8, 97.2}, {66.8, 97.3}, {66.8, 97.3}, {66.8, 97.4}, {66.8, 97.4}, {66.8, 97.5}, {66.8, 97.3}, {66.8, 97.2}, {66.8, 97.1}, {66.8, 97.0}, {66.8, 97.1}, {66.8, 96.9}, {66.8, 96.9}, {66.8, 97.3}, {66.8, 97.3}, {66.8, 97.4}, {66.8, 97.3}, {66.8, 97.5}, {66.8, 97.6}, {66.8, 97.6}, {66.8, 97.5}, {66.8, 97.4}, {66.8, 97.6}, {66.8, 97.8}, {66.8, 97.9}, {66.8, 98.0}, {66.8, 98.0}, {66.8, 97.9}, {66.8, 98.0}, {66.8, 98.0}, {66.8, 98.0}, {66.8, 98.0}, {66.8, 98.0}, {66.8, 98.0}, {66.8, 98.0}, {66.8, 98.1}, {66.8, 98.2}, {66.8, 98.1}, {66.8, 98.1}, {66.8, 98.0}, {66.8, 97.9}, {66.8, 97.9}, {66.8, 97.8}, {66.8, 97.8}, {66.8, 97.9}, {66.8, 97.9}, {66.8, 98.0}, {66.8, 98.1}, {66.8, 98.1}, {66.8, 98.0}, {66.8, 98.0}, {66.8, 97.7}, {66.8, 97.8}, {66.8, 97.9}, {66.8, 97.9}, {66.8, 98.0}, {66.8, 98.1}, {66.8, 98.1}, {66.8, 98.1}, {66.8, 98.1}, {66.8, 72.9, 97.9, 98.2}}, {{15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 60.3}, {15.0, 15.0, 60.3, 60.3}}, {{60.3, 72.9, 72.9, 98.2}, {60.3, 98.2}, {60.3, 98.1}, {60.3, 98.1}, {60.3, 98.3}, {60.3, 98.4}, {60.3, 98.5}, {60.3, 98.4}, {60.3, 98.5}, {60.3, 98.6}, {60.3, 98.6}, {60.3, 98.8}, {60.3, 98.7}, {60.3, 98.7}, {60.3, 98.8}, {60.3, 98.9}, {60.3, 98.6}, {60.3, 98.6}, {60.3, 98.5}, {60.3, 98.4}, {60.3, 98.6}, {60.3, 99.0}, {60.3, 99.0}, {60.3, 98.8}, {60.3, 98.7}, {60.3, 98.6}, {60.3, 98.3}, {60.3, 98.3}, {60.3, 98.4}, {60.3, 98.3}, {60.3, 98.4}, {60.3, 98.4}, {60.3, 98.8}, {60.3, 99.0}, {60.3, 98.8}, {60.3, 98.7}, {60.3, 98.7}, {60.3, 98.5}, {60.3, 98.4}, {60.3, 98.4}, {60.3, 98.5}, {60.3, 98.5}, {60.3, 98.3}, {60.3, 98.4}, {60.3, 99.1}, {60.3, 99.2}, {60.3, 99.3}, {60.3, 99.4}, {60.3, 99.2}, {60.3, 99.0}, {60.3, 99.0}, {60.3, 99.0}, {60.3, 99.0}, {60.3, 98.8}, {60.3, 98.8}, {60.3, 98.8}, {60.3, 98.7}, {60.3, 98.8}, {60.3, 98.9}, {60.3, 98.8}, {60.3, 99.1}, {60.3, 99.1}, {60.3, 99.1}, {60.3, 99.1}, {60.3, 98.9}, {60.3, 98.6}, {60.3, 99.1}, {60.3, 99.0}, {60.3, 98.8}, {60.3, 99.0}, {60.3, 98.9}, {60.3, 98.6}, {60.3, 98.8}, {60.3, 98.8}, {60.3, 98.9}, {60.3, 98.8}, {60.3, 98.5}, {60.3, 98.6}, {60.3, 98.4}, {60.3, 98.4}, {60.3, 98.3}, {60.3, 98.4}, {60.3, 98.3}, {60.3, 98.4}, {60.3, 98.5}, {60.3, 98.5}, {60.3, 98.6}, {60.3, 98.7}, {60.3, 98.6}, {60.3, 98.5}, {60.3, 98.6}, {60.3, 98.6}, {60.3, 98.7}, {60.3, 98.8}, {60.3, 98.9}, {60.3, 99.1}, {60.3, 99.2}, {60.3, 99.1}, {60.3, 99.2}, {60.3, 99.3}, {60.3, 99.3}, {60.3, 99.3}, {60.3, 99.3}, {60.3, 99.2}, {60.3, 99.2}, {60.3, 99.1}, {60.3, 99.2}, {60.3, 99.5}, {60.3, 99.4}, {60.3, 99.4}, {60.3, 99.6}, {60.3, 99.6}, {60.3, 99.6}, {60.3, 99.5}, {60.3, 99.4}, {60.3, 99.3}, {60.3, 99.4}, {60.3, 99.5}, {60.3, 99.5}, {60.3, 99.5}, {60.3, 99.4}, {60.3, 99.6}, {60.3, 99.8}, {60.3, 99.7}, {60.3, 99.7}, {60.3, 99.6}, {60.3, 99.5}, {60.3, 99.8}, {60.3, 99.8}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 99.8}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 99.8}, {60.3, 99.8}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 100.1}, {60.3, 100.0}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 100.0}, {60.3, 99.8}, {60.3, 100.0}, {60.3, 100.1}, {60.3, 100.2}, {60.3, 100.4}, {60.3, 100.4}, {60.3, 100.2}, {60.3, 100.3}, {60.3, 100.4}, {60.3, 100.4}, {60.3, 100.3}, {60.3, 100.3}, {60.3, 100.2}, {60.3, 100.1}, {60.3, 100.1}, {60.3, 99.9}, {60.3, 100.1}, {60.3, 100.0}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 99.7}, {60.3, 99.8}, {60.3, 99.5}, {60.3, 99.6}, {60.3, 99.6}, {60.3, 99.4}, {60.3, 99.7}, {60.3, 99.6}, {60.3, 99.3}, {60.3, 99.3}, {60.3, 99.5}, {60.3, 99.4}, {60.3, 99.3}, {60.3, 99.5}, {60.3, 99.5}, {60.3, 99.5}, {60.3, 99.5}, {60.3, 99.5}, {60.3, 99.4}, {60.3, 99.2}, {60.3, 99.2}, {60.3, 99.3}, {60.3, 99.4}, {60.3, 99.4}, {60.3, 99.5}, {60.3, 99.6}, {60.3, 99.9}, {60.3, 99.8}, {60.3, 99.7}, {60.3, 99.7}, {60.3, 99.7}, {60.3, 99.6}, {60.3, 99.6}, {60.3, 99.7}, {60.3, 99.6}, {60.3, 99.8}, {60.3, 100.0}, {60.3, 100.1}, {60.3, 100.1}, {60.3, 100.2}, {60.3, 100.2}, {60.3, 100.2}, {60.3, 100.3}, {60.3, 100.3}, {60.3, 100.3}, {60.3, 100.2}, {60.3, 100.2}, {60.3, 100.2}, {60.3, 100.2}, {60.3, 100.2}, {60.3, 100.1}, {60.3, 100.0}, {60.3, 99.7}, {60.3, 99.8}, {60.3, 99.9}, {60.3, 99.4}, {60.3, 99.4}, {60.3, 99.9}, {60.3, 100.0}, {60.3, 100.1}, {60.3, 100.2}, {60.3, 100.1}, {60.3, 99.8}, {60.3, 99.1}, {60.3, 98.9}, {60.3, 99.0}, {60.3, 99.3}, {60.3, 99.7}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 100.1}, {60.3, 100.0}, {60.3, 99.8}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 100.2}, {60.3, 100.1}, {60.3, 100.1}, {60.3, 99.8}, {60.3, 99.8}, {60.3, 100.2}, {60.3, 99.9}, {60.3, 100.1}, {60.3, 100.1}, {60.3, 100.2}, {60.3, 100.1}, {60.3, 100.2}, {60.3, 100.0}, {60.3, 100.1}, {60.3, 100.0}, {60.3, 100.2}, {60.3, 100.3}, {60.3, 100.3}, {60.3, 100.3}, {60.3, 100.2}, {60.3, 99.9}, {60.3, 99.9}, {60.3, 100.1}, {60.3, 100.4}, {60.3, 100.5}, {60.3, 100.5}, {60.3, 100.6}, {60.3, 100.5}, {60.3, 100.3}, {60.3, 100.0}, {60.3, 100.0}, {60.3, 100.2}, {60.3, 100.3}, {60.3, 100.6}, {60.3, 100.8}, {60.3, 100.9}, {60.3, 100.9}, {60.3, 100.8}, {60.3, 100.9}, {60.3, 100.6}, {60.3, 100.3}, {60.3, 100.4}, {60.3, 100.9}, {60.3, 101.0}, {60.3, 101.1}, {60.3, 101.1}, {60.3, 101.2}, {60.3, 101.2}, {60.3, 101.3}, {60.3, 101.3}, {60.3, 101.2}, {60.3, 101.1}, {60.3, 101.1}, {60.3, 101.1}, {60.3, 101.1}, {60.3, 101.1}, {60.3, 101.3}, {60.3, 101.4}, {60.3, 101.3}, {60.3, 101.0}, {60.3, 101.2}, {60.3, 101.6}, {60.3, 101.6}, {60.3, 101.6}, {60.3, 101.7}, {60.3, 101.6}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.2}, {60.3, 101.4}, {60.3, 101.3}, {60.3, 101.2}, {60.3, 101.2}, {60.3, 101.4}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.7}, {60.3, 101.8}, {60.3, 101.8}, {60.3, 101.7}, {60.3, 101.8}, {60.3, 101.7}, {60.3, 101.5}, {60.3, 101.4}, {60.3, 101.4}, {60.3, 101.4}, {60.3, 101.4}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.6}, {60.3, 101.6}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.3}, {60.3, 101.2}, {60.3, 101.3}, {60.3, 101.1}, {60.3, 101.0}, {60.3, 101.4}, {60.3, 101.6}, {60.3, 101.5}, {60.3, 101.8}, {60.3, 101.9}, {60.3, 101.9}, {60.3, 101.7}, {60.3, 101.7}, {60.3, 101.7}, {60.3, 101.8}, {60.3, 101.9}, {60.3, 102.0}, {60.3, 102.1}, {60.3, 102.1}, {60.3, 102.1}, {60.3, 101.7}, {60.3, 101.4}, {60.3, 101.3}, {60.3, 101.2}, {60.3, 101.2}, {60.3, 101.1}, {60.3, 100.8}, {60.3, 101.1}, {60.3, 101.2}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.4}, {60.3, 101.3}, {60.3, 101.3}, {60.3, 101.4}, {60.3, 101.7}, {60.3, 101.6}, {60.3, 101.7}, {60.3, 101.5}, {60.3, 101.4}, {60.3, 101.2}, {60.3, 101.2}, {60.3, 101.2}, {60.3, 101.0}, {60.3, 100.9}, {60.3, 100.9}, {60.3, 101.2}, {60.3, 101.3}, {60.3, 101.3}, {60.3, 101.4}, {60.3, 101.6}, {60.3, 101.6}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.4}, {60.3, 101.6}, {60.3, 101.7}, {60.3, 101.8}, {60.3, 101.7}, {60.3, 101.8}, {60.3, 101.7}, {60.3, 101.6}, {60.3, 101.4}, {60.3, 101.7}, {60.3, 101.6}, {60.3, 101.6}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.6}, {60.3, 101.7}, {60.3, 102.0}, {60.3, 102.0}, {60.3, 101.8}, {60.3, 101.9}, {60.3, 101.6}, {60.3, 101.5}, {60.3, 101.5}, {60.3, 101.7}, {60.3, 101.8}, {60.3, 101.7}, {60.3, 101.4}, {60.3, 101.4}, {60.3, 101.7}, {60.3, 102.1}, {60.3, 102.1}, {60.3, 102.0}, {60.3, 102.2}, {60.3, 102.2}, {60.3, 102.3}, {60.3, 102.3}, {60.3, 102.4}, {60.3, 102.3}, {60.3, 102.2}, {60.3, 102.1}, {60.3, 102.2}, {60.3, 102.0}, {60.3, 101.7}, {60.3, 101.8}, {60.3, 102.2}, {60.3, 102.3}, {60.3, 102.0}, {60.3, 102.5}, {60.3, 102.5}, {60.3, 102.3}, {60.3, 102.1}, {60.3, 102.0}, {60.3, 101.8}, {60.3, 101.8}, {60.3, 102.2}, {60.3, 102.4}, {60.3, 102.6}, {60.3, 102.7}, {60.3, 102.9}, {60.3, 102.8}, {60.3, 102.5}, {60.3, 102.3}, {60.3, 102.4}, {60.3, 102.4}, {60.3, 102.2}, {60.3, 102.5}, {60.3, 102.5}, {60.3, 102.6}, {60.3, 102.7}, {60.3, 102.6}, {60.3, 102.4}, {60.3, 102.3}, {60.3, 102.5}, {60.3, 102.4}, {60.3, 102.3}, {60.3, 102.2}, {60.3, 102.0}, {60.3, 102.1}, {60.3, 102.3}, {60.3, 102.2}, {60.3, 102.3}, {60.3, 102.3}, {60.3, 102.4}, {60.3, 102.3}, {60.3, 102.6}, {60.3, 102.7}, {60.3, 102.7}, {60.3, 102.8}, {60.3, 102.7}, {60.3, 102.8}, {60.3, 102.6}, {60.3, 102.7}, {60.3, 102.7}, {60.3, 102.8}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 102.8}, {60.3, 103.1}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.3}, {60.3, 103.2}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.7}, {60.3, 103.7}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.6}, {60.3, 103.6}, {60.3, 103.6}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.3}, {60.3, 103.2}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.0}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 102.8}, {60.3, 102.7}, {60.3, 102.5}, {60.3, 102.4}, {60.3, 102.8}, {60.3, 103.0}, {60.3, 103.1}, {60.3, 103.0}, {60.3, 103.2}, {60.3, 103.1}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.2}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 102.8}, {60.3, 102.9}, {60.3, 103.1}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 102.7}, {60.3, 102.6}, {60.3, 102.6}, {60.3, 102.7}, {60.3, 102.8}, {60.3, 102.8}, {60.3, 102.9}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.2}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 102.6}, {60.3, 102.3}, {60.3, 103.0}, {60.3, 103.1}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 102.9}, {60.3, 102.7}, {60.3, 102.7}, {60.3, 102.7}, {60.3, 102.7}, {60.3, 102.8}, {60.3, 102.9}, {60.3, 102.9}, {60.3, 102.8}, {60.3, 102.8}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 102.9}, {60.3, 102.8}, {60.3, 102.8}, {60.3, 102.8}, {60.3, 103.0}, {60.3, 103.2}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.3}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.2}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.5}, {60.3, 103.8}, {60.3, 103.8}, {60.3, 103.7}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.7}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 104.1}, {60.3, 104.1}, {60.3, 103.9}, {60.3, 103.7}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.7}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 104.0}, {60.3, 104.2}, {60.3, 104.2}, {60.3, 104.1}, {60.3, 104.1}, {60.3, 104.3}, {60.3, 104.4}, {60.3, 104.3}, {60.3, 104.3}, {60.3, 104.3}, {60.3, 104.2}, {60.3, 104.2}, {60.3, 104.1}, {60.3, 104.2}, {60.3, 104.1}, {60.3, 104.1}, {60.3, 104.0}, {60.3, 104.0}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 104.1}, {60.3, 104.1}, {60.3, 104.2}, {60.3, 104.2}, {60.3, 104.3}, {60.3, 104.2}, {60.3, 104.1}, {60.3, 104.0}, {60.3, 104.0}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 104.0}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.7}, {60.3, 103.6}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.7}, {60.3, 103.6}, {60.3, 103.4}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.3}, {60.3, 103.1}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.6}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.7}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 103.7}, {60.3, 103.3}, {60.3, 103.5}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 103.7}, {60.3, 104.1}, {60.3, 104.0}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.6}, {60.3, 103.6}, {60.3, 103.7}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.5}, {60.3, 103.4}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.2}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 102.9}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.2}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.1}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 103.1}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.2}, {60.3, 103.1}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.7}, {60.3, 103.7}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 104.0}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.8}, {60.3, 103.8}, {60.3, 103.7}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 104.0}, {60.3, 104.0}, {60.3, 103.9}, {60.3, 104.1}, {60.3, 104.1}, {60.3, 104.1}, {60.3, 104.2}, {60.3, 104.2}, {60.3, 104.1}, {60.3, 104.1}, {60.3, 104.3}, {60.3, 104.2}, {60.3, 104.3}, {60.3, 104.6}, {60.3, 104.7}, {60.3, 104.7}, {60.3, 104.7}, {60.3, 104.7}, {60.3, 104.7}, {60.3, 104.9}, {60.3, 105.1}, {60.3, 105.2}, {60.3, 105.3}, {60.3, 105.3}, {60.3, 105.3}, {60.3, 105.3}, {60.3, 105.4}, {60.3, 105.5}, {60.3, 105.3}, {60.3, 105.7}, {60.3, 105.8}, {60.3, 105.8}, {60.3, 105.6}, {60.3, 105.7}, {60.3, 105.7}, {60.3, 105.7}, {60.3, 105.7}, {60.3, 105.8}, {60.3, 105.7}, {60.3, 105.5}, {60.3, 105.4}, {60.3, 105.1}, {60.3, 105.2}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.0}, {60.3, 105.0}, {60.3, 104.9}, {60.3, 104.9}, {60.3, 104.7}, {60.3, 104.9}, {60.3, 104.8}, {60.3, 105.0}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.0}, {60.3, 105.0}, {60.3, 105.0}, {60.3, 104.9}, {60.3, 104.9}, {60.3, 104.9}, {60.3, 104.8}, {60.3, 104.8}, {60.3, 104.8}, {60.3, 104.8}, {60.3, 104.7}, {60.3, 104.5}, {60.3, 104.4}, {60.3, 104.2}, {60.3, 104.1}, {60.3, 104.3}, {60.3, 104.4}, {60.3, 104.4}, {60.3, 104.4}, {60.3, 104.3}, {60.3, 104.0}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 103.7}, {60.3, 103.6}, {60.3, 103.5}, {60.3, 103.3}, {60.3, 103.1}, {60.3, 103.1}, {60.3, 103.2}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.1}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 103.0}, {60.3, 102.8}, {60.3, 103.0}, {60.3, 102.9}, {60.3, 103.0}, {60.3, 103.1}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.2}, {60.3, 103.4}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.5}, {60.3, 103.2}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.3}, {60.3, 103.4}, {60.3, 103.4}, {60.3, 103.6}, {60.3, 103.8}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.7}, {60.3, 103.7}, {60.3, 103.8}, {60.3, 103.7}, {60.3, 103.7}, {60.3, 103.8}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 103.8}, {60.3, 103.6}, {60.3, 103.7}, {60.3, 103.8}, {60.3, 103.8}, {60.3, 103.6}, {60.3, 103.8}, {60.3, 104.0}, {60.3, 103.9}, {60.3, 103.9}, {60.3, 104.0}, {60.3, 104.1}, {60.3, 104.2}, {60.3, 104.3}, {60.3, 104.2}, {60.3, 104.2}, {60.3, 104.1}, {60.3, 104.2}, {60.3, 104.3}, {60.3, 104.4}, {60.3, 104.5}, {60.3, 104.2}, {60.3, 104.3}, {60.3, 104.3}, {60.3, 104.7}, {60.3, 104.8}, {60.3, 104.8}, {60.3, 104.8}, {60.3, 104.8}, {60.3, 104.9}, {60.3, 104.8}, {60.3, 104.8}, {60.3, 104.6}, {60.3, 104.5}, {60.3, 104.6}, {60.3, 104.7}, {60.3, 104.9}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 104.9}, {60.3, 104.9}, {60.3, 104.7}, {60.3, 104.7}, {60.3, 104.9}, {60.3, 105.0}, {60.3, 105.0}, {60.3, 105.1}, {60.3, 105.0}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 105.1}, {60.3, 104.9}, {60.3, 105.3}, {60.3, 105.2}, {60.3, 105.3}, {60.3, 105.1}, {60.3, 105.3}, {60.3, 105.2}, {60.3, 105.3}, {60.3, 105.2}, {60.3, 105.3}, {60.3, 105.4}, {60.3, 105.4}, {60.3, 105.5}, {60.3, 105.6}, {60.3, 105.5}, {60.3, 105.5}, {60.3, 105.3}, {60.3, 105.4}, {60.3, 105.4}, {60.3, 105.5}, {60.3, 105.5}, {60.3, 105.6}, {60.3, 105.6}, {60.3, 105.6}, {60.3, 105.6}, {60.3, 105.6}, {60.3, 105.5}, {60.3, 105.6}, {60.3, 105.6}, {60.3, 105.6}, {60.3, 105.5}, {60.3, 105.7}, {60.3, 105.9}, {60.3, 105.9}, {60.3, 106.0}, {60.3, 106.0}, {60.3, 106.0}, {60.3, 106.0}, {60.3, 105.9}, {60.3, 105.9}, {60.3, 106.0}, {60.3, 106.2}, {60.3, 106.5}, {60.3, 106.5}, {60.3, 106.4}, {60.3, 106.4}, {60.3, 106.3}, {60.3, 106.2}, {60.3, 106.1}, {60.3, 106.3}, {60.3, 106.3}, {60.3, 106.2}, {60.3, 106.3}, {60.3, 106.3}, {60.3, 106.3}, {60.3, 106.3}, {60.3, 106.3}, {60.3, 106.3}, {60.3, 106.4}, {60.3, 106.4}, {60.3, 106.4}, {60.3, 106.3}, {60.3, 106.0}, {60.3, 106.5}, {60.3, 106.5}, {60.3, 106.4}, {60.3, 106.4}, {60.3, 106.6}, {60.3, 106.8}, {60.3, 106.8}, {60.3, 106.7}, {60.3, 106.6}, {60.3, 106.7}, {60.3, 106.7}, {60.3, 106.6}, {60.3, 106.6}, {60.3, 106.7}, {60.3, 106.7}, {60.3, 106.7}, {60.3, 106.9}, {60.3, 106.7}, {60.3, 106.5}, {60.3, 106.8}, {60.3, 107.0}, {60.3, 107.0}, {60.3, 107.1}, {60.3, 107.1}, {60.3, 107.2}, {60.3, 107.0}, {60.3, 106.8}, {60.3, 106.7}, {60.3, 107.1}, {60.3, 106.9}, {60.3, 106.8}, {60.3, 106.8}, {60.3, 106.8}, {60.3, 107.2}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.4}, {60.3, 107.3}, {60.3, 107.2}, {60.3, 107.1}, {60.3, 107.1}, {60.3, 107.1}, {60.3, 107.1}, {60.3, 107.1}, {60.3, 107.1}, {60.3, 107.2}, {60.3, 107.2}, {60.3, 107.1}, {60.3, 107.0}, {60.3, 107.0}, {60.3, 107.2}, {60.3, 107.3}, {60.3, 107.3}, {60.3, 107.3}, {60.3, 107.4}, {60.3, 107.3}, {60.3, 107.3}, {60.3, 107.3}, {60.3, 107.2}, {60.3, 107.3}, {60.3, 107.4}, {60.3, 107.3}, {60.3, 107.3}, {60.3, 107.6}, {60.3, 107.7}, {60.3, 107.8}, {60.3, 107.8}, {60.3, 107.7}, {60.3, 107.6}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.6}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.6}, {60.3, 107.6}, {60.3, 107.5}, {60.3, 107.6}, {60.3, 107.5}, {60.3, 107.6}, {60.3, 107.6}, {60.3, 107.6}, {60.3, 107.5}, {60.3, 107.4}, {60.3, 107.4}, {60.3, 107.4}, {60.3, 107.4}, {60.3, 107.4}, {60.3, 107.3}, {60.3, 107.1}, {60.3, 107.1}, {60.3, 107.0}, {60.3, 107.2}, {60.3, 107.3}, {60.3, 107.4}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.6}, {60.3, 107.5}, {60.3, 107.3}, {60.3, 107.3}, {60.3, 107.5}, {60.3, 107.4}, {60.3, 107.4}, {60.3, 107.3}, {60.3, 107.4}, {60.3, 107.6}, {60.3, 107.5}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.6}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.6}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.8}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.8}, {60.3, 107.8}, {60.3, 107.6}, {60.3, 107.6}, {60.3, 107.8}, {60.3, 108.0}, {60.3, 108.0}, {60.3, 108.0}, {60.3, 108.0}, {60.3, 107.9}, {60.3, 107.8}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.8}, {60.3, 107.7}, {60.3, 107.6}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.5}, {60.3, 107.6}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.7}, {60.3, 107.8}, {60.3, 107.9}, {60.3, 107.9}, {60.3, 107.9}, {60.3, 108.0}, {60.3, 107.9}, {60.3, 107.9}, {60.3, 107.8}, {60.3, 107.6}, {60.3, 107.6}, {60.3, 107.6}, {60.3, 107.7}, {60.3, 107.9}, {60.3, 108.0}, {60.3, 108.2}, {60.3, 108.4}, {60.3, 108.5}, {60.3, 108.6}, {60.3, 108.5}, {60.3, 108.5}, {60.3, 108.6}, {60.3, 108.5}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.9}, {60.3, 108.9}, {60.3, 108.7}, {60.3, 108.7}, {60.3, 108.6}, {60.3, 108.7}, {60.3, 108.6}, {60.3, 108.5}, {60.3, 108.5}, {60.3, 108.3}, {60.3, 108.3}, {60.3, 108.4}, {60.3, 108.3}, {60.3, 108.4}, {60.3, 108.4}, {60.3, 108.4}, {60.3, 108.4}, {60.3, 108.4}, {60.3, 108.4}, {60.3, 108.4}, {60.3, 108.4}, {60.3, 108.3}, {60.3, 108.2}, {60.3, 108.1}, {60.3, 108.3}, {60.3, 108.5}, {60.3, 108.5}, {60.3, 108.5}, {60.3, 108.4}, {60.3, 108.6}, {60.3, 108.5}, {60.3, 108.6}, {60.3, 108.6}, {60.3, 108.7}, {60.3, 108.8}, {60.3, 109.0}, {60.3, 109.0}, {60.3, 108.9}, {60.3, 108.8}, {60.3, 108.7}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.7}, {60.3, 108.6}, {60.3, 108.6}, {60.3, 108.6}, {60.3, 108.8}, {60.3, 108.6}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.7}, {60.3, 108.6}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.9}, {60.3, 109.0}, {60.3, 109.0}, {60.3, 109.0}, {60.3, 108.9}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.8}, {60.3, 108.9}, {60.3, 109.1}, {60.3, 109.3}, {60.3, 109.3}, {60.3, 109.5}, {60.3, 109.6}, {60.3, 109.5}, {60.3, 109.4}, {60.3, 109.5}, {60.3, 109.5}, {60.3, 109.3}, {60.3, 109.3}, {60.3, 109.3}, {60.3, 109.5}, {60.3, 109.5}, {60.3, 109.4}, {60.3, 109.5}, {60.3, 109.5}, {60.3, 109.4}, {60.3, 109.3}, {60.3, 109.1}, {60.3, 109.2}, {60.3, 109.2}, {60.3, 109.1}, {60.3, 109.1}, {60.3, 109.0}, {60.3, 108.8}, {60.3, 108.6}, {60.3, 108.7}, {60.3, 108.7}, {60.3, 108.8}, {60.3, 108.9}, {60.3, 108.9}, {60.3, 109.0}, {60.3, 108.9}, {60.3, 108.9}, {60.3, 108.9}, {60.3, 108.9}, {60.3, 109.0}, {60.3, 109.0}, {60.3, 109.1}, {60.3, 109.1}, {60.3, 109.1}, {60.3, 109.1}, {60.3, 108.9}, {60.3, 108.8}, {60.3, 108.6}, {60.3, 108.7}, {60.3, 108.9}, {60.3, 109.0}, {60.3, 109.0}, {60.3, 109.1}, {60.3, 109.1}, {60.3, 109.0}, {60.3, 109.2}, {60.3, 109.2}, {60.3, 109.3}, {60.3, 109.4}, {60.3, 109.3}, {60.3, 109.3}, {60.3, 109.3}, {60.3, 109.3}, {60.3, 109.4}, {60.3, 109.4}, {60.3, 109.5}, {60.3, 109.6}, {60.3, 109.7}, {60.3, 109.8}, {60.3, 109.6}, {60.3, 109.5}, {60.3, 109.3}, {60.3, 109.4}, {60.3, 109.6}, {60.3, 109.9}, {60.3, 110.0}, {60.3, 110.1}, {60.3, 110.2}, {60.3, 110.2}, {60.3, 110.2}, {60.3, 110.3}, {60.3, 110.1}, {60.3, 110.2}, {60.3, 110.4}, {60.3, 110.5}, {60.3, 110.8}, {60.3, 110.9}, {60.3, 110.9}, {60.3, 111.1}, {60.3, 111.1}, {60.3, 111.3}, {60.3, 111.2}, {60.3, 111.2}, {60.3, 111.2}, {60.3, 111.4}, {60.3, 111.5}, {60.3, 111.4}, {60.3, 111.2}, {60.3, 110.6}, {60.3, 110.5}, {60.3, 111.1}, {60.3, 111.2}, {60.3, 111.2}, {60.3, 111.3}, {60.3, 111.3}, {60.3, 111.5}, {60.3, 111.5}, {60.3, 111.4}, {60.3, 111.5}, {60.3, 111.5}, {60.3, 111.5}, {60.3, 111.4}, {60.3, 111.2}, {60.3, 111.2}, {60.3, 111.3}, {60.3, 111.4}, {60.3, 111.6}, {60.3, 111.4}, {60.3, 111.8}, {60.3, 112.0}, {60.3, 112.1}, {60.3, 112.2}, {60.3, 112.1}, {60.3, 112.2}, {60.3, 112.3}, {60.3, 112.4}, {60.3, 112.4}, {60.3, 112.5}, {60.3, 112.4}, {60.3, 112.4}, {60.3, 112.8}, {60.3, 112.7}, {60.3, 112.7}, {60.3, 112.8}, {60.3, 112.8}, {60.3, 112.9}, {60.3, 112.7}, {60.3, 112.7}, {60.3, 112.6}, {60.3, 112.6}, {60.3, 112.5}, {60.3, 112.6}, {60.3, 112.5}, {60.3, 112.6}, {60.3, 112.6}, {60.3, 112.6}, {60.3, 112.7}, {60.3, 112.8}, {60.3, 112.8}, {60.3, 112.8}, {60.3, 112.9}, {60.3, 113.0}, {60.3, 112.9}, {60.3, 112.5}, {60.3, 112.5}, {60.3, 112.5}, {60.3, 112.6}, {60.3, 112.6}, {60.3, 112.7}, {60.3, 113.0}, {60.3, 113.2}, {60.3, 113.2}, {60.3, 113.3}, {60.3, 113.3}, {60.3, 113.4}, {60.3, 113.5}, {60.3, 113.5}, {60.3, 113.5}, {60.3, 113.7}, {60.3, 113.8}, {60.3, 113.8}, {60.3, 113.8}, {60.3, 113.8}, {60.3, 114.1}, {60.3, 114.1}, {60.3, 114.1}, {60.3, 114.1}, {60.3, 114.3}, {60.3, 114.6}, {60.3, 114.5}, {60.3, 114.6}, {60.3, 114.6}, {60.3, 114.7}, {60.3, 114.6}, {60.3, 114.7}, {60.3, 114.6}, {60.3, 114.7}, {60.3, 114.5}, {60.3, 114.5}, {60.3, 114.5}, {60.3, 114.5}, {60.3, 114.5}, {60.3, 114.5}, {60.3, 114.4}, {60.3, 114.3}, {60.3, 114.4}, {60.3, 114.7}, {60.3, 114.9}, {60.3, 115.0}, {60.3, 115.2}, {60.3, 115.2}, {60.3, 115.4}, {60.3, 115.2}, {60.3, 115.1}, {60.3, 115.1}, {60.3, 115.3}, {60.3, 115.4}, {60.3, 115.5}, {60.3, 115.7}, {60.3, 115.7}, {60.3, 115.8}, {60.3, 115.9}, {60.3, 115.9}, {60.3, 115.8}, {60.3, 115.8}, {60.3, 115.8}, {60.3, 115.8}, {60.3, 115.9}, {60.3, 115.8}, {60.3, 115.8}, {60.3, 115.7}, {60.3, 115.6}, {60.3, 115.6}, {60.3, 115.8}, {60.3, 115.8}, {60.3, 115.8}, {60.3, 115.7}, {60.3, 115.7}, {60.3, 115.6}, {60.3, 115.6}, {60.3, 115.6}, {60.3, 115.6}, {60.3, 115.7}, {60.3, 115.8}, {60.3,  60.3, 115.9, 115.9}};
		}
	}
}
