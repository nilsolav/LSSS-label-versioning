netcdf mask {
	:date_created = "20190819T134900Z";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200728T132547";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 3;
			channels = 4;
			categories = 12;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  12.0, 12.0, 76.9;
			max_depth =  91.7, 102.0,  85.1;
			start_time = 128216212101214208, 128216192551214208, 128216215781214208;
			end_time = 128216226481214208, 128216212101214208, 128216215821214208;
			region_id = 1, 2, 3;
			region_name = "Layer1","Layer2","Layer1";
			region_provenance = "LSSS", "LSSS", "LSSS";
			region_comment = "", "", "";
			region_category_names = "0", "0", "0", "0", "0", "0", "0", "0", "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1,  2,  3,  4,  5,  6,  7,  8,  9, 10, 11, 12;
			region_type = analysis, analysis, analysis;
			channel_names = "18", "38", "120", "200";
			region_channels = 15, 15, 15;
			mask_times = {1.282162121012142e+17, 1.282162121112142e+17, 1.282162121212143e+17, 1.282162121312142e+17, 1.282162121412142e+17, 1.282162121512142e+17, 1.282162121612143e+17, 1.282162121712142e+17, 1.282162121812143e+17, 1.282162121912142e+17, 1.282162122012143e+17, 1.282162122112142e+17, 1.282162122212142e+17, 1.282162122312143e+17, 1.282162122412142e+17, 1.282162122512142e+17, 1.282162122612142e+17, 1.282162122712143e+17, 1.282162122812142e+17, 1.282162122912143e+17, 1.282162123012142e+17, 1.282162123112143e+17, 1.282162123212142e+17, 1.282162123312143e+17, 1.282162123412142e+17, 1.282162123512142e+17, 1.282162123612142e+17, 1.282162123712142e+17, 1.282162123812143e+17, 1.282162123912142e+17, 1.282162124012142e+17, 1.282162124112142e+17, 1.282162124212143e+17, 1.282162124312142e+17, 1.282162124412143e+17, 1.282162124512142e+17, 1.282162124612143e+17, 1.282162124712142e+17, 1.282162124812142e+17, 1.282162124912143e+17, 1.282162125012142e+17, 1.282162125112142e+17, 1.282162125212142e+17, 1.282162125312143e+17, 1.282162125412142e+17, 1.282162125512143e+17, 1.282162125612142e+17, 1.282162125712143e+17, 1.282162125812142e+17, 1.282162125912143e+17, 1.282162126012142e+17, 1.282162126112142e+17, 1.282162126212142e+17, 1.282162126312142e+17, 1.282162126412143e+17, 1.282162126512142e+17, 1.282162126612142e+17, 1.282162126712142e+17, 1.282162126812143e+17, 1.282162126912142e+17, 1.282162127012143e+17, 1.282162127112142e+17, 1.282162127212143e+17, 1.282162127312142e+17, 1.282162127412142e+17, 1.282162127512143e+17, 1.282162127612142e+17, 1.282162127712142e+17, 1.282162127812142e+17, 1.282162127912143e+17, 1.282162128012142e+17, 1.282162128112143e+17, 1.282162128212142e+17, 1.282162128312143e+17, 1.282162128412142e+17, 1.282162128512142e+17, 1.282162128612143e+17, 1.282162128712142e+17, 1.282162128812142e+17, 1.282162128912142e+17, 1.282162129012143e+17, 1.282162129112142e+17, 1.282162129212143e+17, 1.282162129312142e+17, 1.282162129412143e+17, 1.282162129512142e+17, 1.282162129612143e+17, 1.282162129712142e+17, 1.282162129812142e+17, 1.282162129912142e+17, 1.282162130012142e+17, 1.282162130112143e+17, 1.282162130212142e+17, 1.282162130312142e+17, 1.282162130412142e+17, 1.282162130512143e+17, 1.282162130612142e+17, 1.282162130712143e+17, 1.282162130812142e+17, 1.282162130912143e+17, 1.282162131012142e+17, 1.282162131112142e+17, 1.282162131212143e+17, 1.282162131312142e+17, 1.282162131412142e+17, 1.282162131512142e+17, 1.282162131612143e+17, 1.282162131712142e+17, 1.282162131812143e+17, 1.282162131912142e+17, 1.282162132012143e+17, 1.282162132112142e+17, 1.282162132212143e+17, 1.282162132312142e+17, 1.282162132412142e+17, 1.282162132512142e+17, 1.282162132612142e+17, 1.282162132712143e+17, 1.282162132812142e+17, 1.282162132912142e+17, 1.282162133012142e+17, 1.282162133112143e+17, 1.282162133212142e+17, 1.282162133312143e+17, 1.282162133412142e+17, 1.282162133512143e+17, 1.282162133612142e+17, 1.282162133712142e+17, 1.282162133812143e+17, 1.282162133912142e+17, 1.282162134012142e+17, 1.282162134112142e+17, 1.282162134212143e+17, 1.282162134312142e+17, 1.282162134412143e+17, 1.282162134512142e+17, 1.282162134612143e+17, 1.282162134712142e+17, 1.282162134812143e+17, 1.282162134912142e+17, 1.282162135012142e+17, 1.282162135112142e+17, 1.282162135212142e+17, 1.282162135312143e+17, 1.282162135412142e+17, 1.282162135512142e+17, 1.282162135612142e+17, 1.282162135712143e+17, 1.282162135812142e+17, 1.282162135912143e+17, 1.282162136012142e+17, 1.282162136112143e+17, 1.282162136212142e+17, 1.282162136312142e+17, 1.282162136412143e+17, 1.282162136512142e+17, 1.282162136612142e+17, 1.282162136712142e+17, 1.282162136812143e+17, 1.282162136912142e+17, 1.282162137012143e+17, 1.282162137112142e+17, 1.282162137212143e+17, 1.282162137312142e+17, 1.282162137412142e+17, 1.282162137512143e+17, 1.282162137612142e+17, 1.282162137712142e+17, 1.282162137812142e+17, 1.282162137912143e+17, 1.282162138012142e+17, 1.282162138112142e+17, 1.282162138212142e+17, 1.282162138312143e+17, 1.282162138412142e+17, 1.282162138512143e+17, 1.282162138612142e+17, 1.282162138712142e+17, 1.282162138812142e+17, 1.282162138912142e+17, 1.282162139012143e+17, 1.282162139112142e+17, 1.282162139212142e+17, 1.282162139312142e+17, 1.282162139412143e+17, 1.282162139512142e+17, 1.282162139612143e+17, 1.282162139712142e+17, 1.282162139812143e+17, 1.282162139912142e+17, 1.282162140012142e+17, 1.282162140112143e+17, 1.282162140212142e+17, 1.282162140312142e+17, 1.282162140412142e+17, 1.282162140512143e+17, 1.282162140612142e+17, 1.282162140712143e+17, 1.282162140812142e+17, 1.282162140912143e+17, 1.282162141012142e+17, 1.282162141112143e+17, 1.282162141212142e+17, 1.282162141312142e+17, 1.282162141412142e+17, 1.282162141512142e+17, 1.282162141612143e+17, 1.282162141712142e+17, 1.282162141812142e+17, 1.282162141912142e+17, 1.282162142012143e+17, 1.282162142112142e+17, 1.282162142212143e+17, 1.282162142312142e+17, 1.282162142412143e+17, 1.282162142512142e+17, 1.282162142612142e+17, 1.282162142712143e+17, 1.282162142812142e+17, 1.282162142912142e+17, 1.282162143012142e+17, 1.282162143112143e+17, 1.282162143212142e+17, 1.282162143312143e+17, 1.282162143412142e+17, 1.282162143512143e+17, 1.282162143612142e+17, 1.282162143712143e+17, 1.282162143812142e+17, 1.282162143912142e+17, 1.282162144012142e+17, 1.282162144112142e+17, 1.282162144212143e+17, 1.282162144312142e+17, 1.282162144412142e+17, 1.282162144512142e+17, 1.282162144612143e+17, 1.282162144712142e+17, 1.282162144812143e+17, 1.282162144912142e+17, 1.282162145012143e+17, 1.282162145112142e+17, 1.282162145212142e+17, 1.282162145312143e+17, 1.282162145412142e+17, 1.282162145512142e+17, 1.282162145612142e+17, 1.282162145712143e+17, 1.282162145812142e+17, 1.282162145912143e+17, 1.282162146012142e+17, 1.282162146112143e+17, 1.282162146212142e+17, 1.282162146312143e+17, 1.282162146412143e+17, 1.282162146512142e+17, 1.282162146612142e+17, 1.282162146712142e+17, 1.282162146812143e+17, 1.282162146912142e+17, 1.282162147012142e+17, 1.282162147112142e+17, 1.282162147212143e+17, 1.282162147312142e+17, 1.282162147412143e+17, 1.282162147512142e+17, 1.282162147612142e+17, 1.282162147712142e+17, 1.282162147812142e+17, 1.282162147912143e+17, 1.282162148012142e+17, 1.282162148112142e+17, 1.282162148212142e+17, 1.282162148312143e+17, 1.282162148412142e+17, 1.282162148512143e+17, 1.282162148612142e+17, 1.282162148712143e+17, 1.282162148812142e+17, 1.282162148912142e+17, 1.282162149012143e+17, 1.282162149112142e+17, 1.282162149212142e+17, 1.282162149312142e+17, 1.282162149412143e+17, 1.282162149512142e+17, 1.282162149612143e+17, 1.282162149712142e+17, 1.282162149812143e+17, 1.282162149912142e+17, 1.282162150012143e+17, 1.282162150112142e+17, 1.282162150212142e+17, 1.282162150312142e+17, 1.282162150412142e+17, 1.282162150512143e+17, 1.282162150612142e+17, 1.282162150712142e+17, 1.282162150812142e+17, 1.282162150912143e+17, 1.282162151012142e+17, 1.282162151112143e+17, 1.282162151212142e+17, 1.282162151312143e+17, 1.282162151412142e+17, 1.282162151512142e+17, 1.282162151612143e+17, 1.282162151712142e+17, 1.282162151812142e+17, 1.282162151912142e+17, 1.282162152012143e+17, 1.282162152112142e+17, 1.282162152212143e+17, 1.282162152312142e+17, 1.282162152412143e+17, 1.282162152512142e+17, 1.282162152612143e+17, 1.282162152712142e+17, 1.282162152812142e+17, 1.282162152912142e+17, 1.282162153012142e+17, 1.282162153112143e+17, 1.282162153212142e+17, 1.282162153312142e+17, 1.282162153412142e+17, 1.282162153512143e+17, 1.282162153612142e+17, 1.282162153712143e+17, 1.282162153812142e+17, 1.282162153912143e+17, 1.282162154012142e+17, 1.282162154112142e+17, 1.282162154212143e+17, 1.282162154312142e+17, 1.282162154412142e+17, 1.282162154512142e+17, 1.282162154612143e+17, 1.282162154712142e+17, 1.282162154812143e+17, 1.282162154912142e+17, 1.282162155012143e+17, 1.282162155112142e+17, 1.282162155212143e+17, 1.282162155312142e+17, 1.282162155412142e+17, 1.282162155512142e+17, 1.282162155612142e+17, 1.282162155712143e+17, 1.282162155812142e+17, 1.282162155912142e+17, 1.282162156012142e+17, 1.282162156112143e+17, 1.282162156212142e+17, 1.282162156312143e+17, 1.282162156412142e+17, 1.282162156512142e+17, 1.282162156612142e+17, 1.282162156712142e+17, 1.282162156812143e+17, 1.282162156912142e+17, 1.282162157012142e+17, 1.282162157112142e+17, 1.282162157212143e+17, 1.282162157312142e+17, 1.282162157512142e+17, 1.282162157612143e+17, 1.282162157712142e+17, 1.282162157812142e+17, 1.282162157912143e+17, 1.282162158012142e+17, 1.282162158112142e+17, 1.282162158212142e+17, 1.282162158312143e+17, 1.282162158412142e+17, 1.282162158512143e+17, 1.282162158612142e+17, 1.282162158712143e+17, 1.282162158812142e+17, 1.282162158912143e+17, 1.282162159012142e+17, 1.282162159112142e+17, 1.282162159212142e+17, 1.282162159312142e+17, 1.282162159412143e+17, 1.282162159512142e+17, 1.282162159612142e+17, 1.282162159712142e+17, 1.282162159812143e+17, 1.282162159912142e+17, 1.282162160012143e+17, 1.282162160112142e+17, 1.282162160212143e+17, 1.282162160312142e+17, 1.282162160412142e+17, 1.282162160512143e+17, 1.282162160612142e+17, 1.282162160712142e+17, 1.282162160812142e+17, 1.282162160912143e+17, 1.282162161012142e+17, 1.282162161112143e+17, 1.282162161212142e+17, 1.282162161312143e+17, 1.282162161412142e+17, 1.282162161512143e+17, 1.282162161612142e+17, 1.282162161712142e+17, 1.282162161812142e+17, 1.282162161912142e+17, 1.282162162012143e+17, 1.282162162112142e+17, 1.282162162212142e+17, 1.282162162312142e+17, 1.282162162412143e+17, 1.282162162512142e+17, 1.282162162612143e+17, 1.282162162712142e+17, 1.282162162812143e+17, 1.282162162912142e+17, 1.282162163012142e+17, 1.282162163112143e+17, 1.282162163212142e+17, 1.282162163312142e+17, 1.282162163412142e+17, 1.282162163512143e+17, 1.282162163612142e+17, 1.282162163712143e+17, 1.282162163812142e+17, 1.282162163912143e+17, 1.282162164012142e+17, 1.282162164112143e+17, 1.282162164212142e+17, 1.282162164312142e+17, 1.282162164412142e+17, 1.282162164512142e+17, 1.282162164612143e+17, 1.282162164712142e+17, 1.282162164812142e+17, 1.282162164912142e+17, 1.282162165012143e+17, 1.282162165112142e+17, 1.282162165212143e+17, 1.282162165312142e+17, 1.282162165412143e+17, 1.282162165512142e+17, 1.282162165612142e+17, 1.282162165712143e+17, 1.282162165812142e+17, 1.282162165912142e+17, 1.282162166012142e+17, 1.282162166112143e+17, 1.282162166212142e+17, 1.282162166312143e+17, 1.282162166412142e+17, 1.282162166512143e+17, 1.282162166612142e+17, 1.282162166712142e+17, 1.282162166812143e+17, 1.282162166912142e+17, 1.282162167012142e+17, 1.282162167112142e+17, 1.282162167212143e+17, 1.282162167312142e+17, 1.282162167412143e+17, 1.282162167512142e+17, 1.282162167612143e+17, 1.282162167712142e+17, 1.282162167812143e+17, 1.282162167912142e+17, 1.282162168012142e+17, 1.282162168112142e+17, 1.282162168212142e+17, 1.282162168312143e+17, 1.282162168412142e+17, 1.282162168512142e+17, 1.282162168612142e+17, 1.282162168712143e+17, 1.282162168812142e+17, 1.282162168912143e+17, 1.282162169012142e+17, 1.282162169112143e+17, 1.282162169212142e+17, 1.282162169312142e+17, 1.282162169412143e+17, 1.282162169512142e+17, 1.282162169612142e+17, 1.282162169712142e+17, 1.282162169812143e+17, 1.282162169912142e+17, 1.282162170012143e+17, 1.282162170112142e+17, 1.282162170212143e+17, 1.282162170312142e+17, 1.282162170412143e+17, 1.282162170512142e+17, 1.282162170612142e+17, 1.282162170712142e+17, 1.282162170812142e+17, 1.282162170912143e+17, 1.282162171012142e+17, 1.282162171112142e+17, 1.282162171212142e+17, 1.282162171312143e+17, 1.282162171412142e+17, 1.282162171512143e+17, 1.282162171612142e+17, 1.282162171712143e+17, 1.282162171812142e+17, 1.282162171912142e+17, 1.282162172012143e+17, 1.282162172112142e+17, 1.282162172212142e+17, 1.282162172312142e+17, 1.282162172412143e+17, 1.282162172512142e+17, 1.282162172612143e+17, 1.282162172712142e+17, 1.282162172812143e+17, 1.282162172912142e+17, 1.282162173012143e+17, 1.282162173112142e+17, 1.282162173212142e+17, 1.282162173312142e+17, 1.282162173412142e+17, 1.282162173512143e+17, 1.282162173612142e+17, 1.282162173712142e+17, 1.282162173812142e+17, 1.282162173912143e+17, 1.282162174012142e+17, 1.282162174112143e+17, 1.282162174212142e+17, 1.282162174312143e+17, 1.282162174412142e+17, 1.282162174512142e+17, 1.282162174612143e+17, 1.282162174712142e+17, 1.282162174812142e+17, 1.282162174912142e+17, 1.282162175012143e+17, 1.282162175112142e+17, 1.282162175212143e+17, 1.282162175312142e+17, 1.282162175412143e+17, 1.282162175512142e+17, 1.282162175612142e+17, 1.282162175712143e+17, 1.282162175812142e+17, 1.282162175912142e+17, 1.282162176012142e+17, 1.282162176112143e+17, 1.282162176212142e+17, 1.282162176312142e+17, 1.282162176412142e+17, 1.282162176512143e+17, 1.282162176612142e+17, 1.282162176712143e+17, 1.282162176812142e+17, 1.282162176912142e+17, 1.282162177012142e+17, 1.282162177112142e+17, 1.282162177212143e+17, 1.282162177312142e+17, 1.282162177412142e+17, 1.282162177512142e+17, 1.282162177612143e+17, 1.282162177712142e+17, 1.282162177812143e+17, 1.282162177912142e+17, 1.282162178012143e+17, 1.282162178112142e+17, 1.282162178212142e+17, 1.282162178312143e+17, 1.282162178412142e+17, 1.282162178512142e+17, 1.282162178612142e+17, 1.282162178712143e+17, 1.282162178812142e+17, 1.282162178912143e+17, 1.282162179012142e+17, 1.282162179112143e+17, 1.282162179212142e+17, 1.282162179312143e+17, 1.282162179412142e+17, 1.282162179512142e+17, 1.282162179612142e+17, 1.282162179712142e+17, 1.282162179812143e+17, 1.282162179912142e+17, 1.282162180012142e+17, 1.282162180112142e+17, 1.282162180212143e+17, 1.282162180312142e+17, 1.282162180412143e+17, 1.282162180512142e+17, 1.282162180612143e+17, 1.282162180712142e+17, 1.282162180812142e+17, 1.282162180912143e+17, 1.282162181012142e+17, 1.282162181112142e+17, 1.282162181212142e+17, 1.282162181312143e+17, 1.282162181412142e+17, 1.282162181512143e+17, 1.282162181612142e+17, 1.282162181712143e+17, 1.282162181812142e+17, 1.282162181912143e+17, 1.282162182012142e+17, 1.282162182112142e+17, 1.282162182212142e+17, 1.282162182312142e+17, 1.282162182412143e+17, 1.282162182512142e+17, 1.282162182612142e+17, 1.282162182712142e+17, 1.282162182812143e+17, 1.282162182912142e+17, 1.282162183012143e+17, 1.282162183112142e+17, 1.282162183212143e+17, 1.282162183312142e+17, 1.282162183412142e+17, 1.282162183512143e+17, 1.282162183612142e+17, 1.282162183712142e+17, 1.282162183812142e+17, 1.282162183912143e+17, 1.282162184012142e+17, 1.282162184112143e+17, 1.282162184212142e+17, 1.282162184312143e+17, 1.282162184412142e+17, 1.282162184512143e+17, 1.282162184612143e+17, 1.282162184712142e+17, 1.282162184812142e+17, 1.282162184912142e+17, 1.282162185012143e+17, 1.282162185112142e+17, 1.282162185212142e+17, 1.282162185312142e+17, 1.282162185412143e+17, 1.282162185512142e+17, 1.282162185612143e+17, 1.282162185712142e+17, 1.282162185812142e+17, 1.282162185912142e+17, 1.282162186012142e+17, 1.282162186112143e+17, 1.282162186212142e+17, 1.282162186312142e+17, 1.282162186412142e+17, 1.282162186512143e+17, 1.282162186612142e+17, 1.282162186712143e+17, 1.282162186812142e+17, 1.282162186912143e+17, 1.282162187012142e+17, 1.282162187112142e+17, 1.282162187212143e+17, 1.282162187312142e+17, 1.282162187412142e+17, 1.282162187512142e+17, 1.282162187612143e+17, 1.282162187712142e+17, 1.282162187812143e+17, 1.282162187912142e+17, 1.282162188012143e+17, 1.282162188112142e+17, 1.282162188212143e+17, 1.282162188312142e+17, 1.282162188412142e+17, 1.282162188512142e+17, 1.282162188612142e+17, 1.282162188712143e+17, 1.282162188812142e+17, 1.282162188912142e+17, 1.282162189012142e+17, 1.282162189112143e+17, 1.282162189212142e+17, 1.282162189312143e+17, 1.282162189412142e+17, 1.282162189512143e+17, 1.282162189612142e+17, 1.282162189712142e+17, 1.282162189812143e+17, 1.282162189912142e+17, 1.282162190012142e+17, 1.282162190112142e+17, 1.282162190212143e+17, 1.282162190312142e+17, 1.282162190412143e+17, 1.282162190512142e+17, 1.282162190612143e+17, 1.282162190712142e+17, 1.282162190812143e+17, 1.282162190912142e+17, 1.282162191012142e+17, 1.282162191112142e+17, 1.282162191212142e+17, 1.282162191312143e+17, 1.282162191412142e+17, 1.282162191512142e+17, 1.282162191612142e+17, 1.282162191712143e+17, 1.282162191812142e+17, 1.282162191912143e+17, 1.282162192012142e+17, 1.282162192112143e+17, 1.282162192212142e+17, 1.282162192312142e+17, 1.282162192412143e+17, 1.282162192512142e+17, 1.282162192612142e+17, 1.282162192712142e+17, 1.282162192812143e+17, 1.282162192912142e+17, 1.282162193012143e+17, 1.282162193112142e+17, 1.282162193212143e+17, 1.282162193312142e+17, 1.282162193412143e+17, 1.282162193512142e+17, 1.282162193612142e+17, 1.282162193712142e+17, 1.282162193812142e+17, 1.282162193912143e+17, 1.282162194012142e+17, 1.282162194112142e+17, 1.282162194212142e+17, 1.282162194312143e+17, 1.282162194412142e+17, 1.282162194512143e+17, 1.282162194612142e+17, 1.282162194712143e+17, 1.282162194812142e+17, 1.282162194912142e+17, 1.282162195012143e+17, 1.282162195112142e+17, 1.282162195212142e+17, 1.282162195312142e+17, 1.282162195412143e+17, 1.282162195512142e+17, 1.282162195612143e+17, 1.282162195712142e+17, 1.282162195812143e+17, 1.282162195912142e+17, 1.282162196012142e+17, 1.282162196112143e+17, 1.282162196212142e+17, 1.282162196312142e+17, 1.282162196412142e+17, 1.282162196512143e+17, 1.282162196612142e+17, 1.282162196712143e+17, 1.282162196812142e+17, 1.282162196912143e+17, 1.282162197012142e+17, 1.282162197112143e+17, 1.282162197212142e+17, 1.282162197312142e+17, 1.282162197412142e+17, 1.282162197512142e+17, 1.282162197612143e+17, 1.282162197712142e+17, 1.282162197812142e+17, 1.282162197912142e+17, 1.282162198012143e+17, 1.282162198112142e+17, 1.282162198212143e+17, 1.282162198312142e+17, 1.282162198412143e+17, 1.282162198512142e+17, 1.282162198612142e+17, 1.282162198712143e+17, 1.282162198812142e+17, 1.282162198912142e+17, 1.282162199012142e+17, 1.282162199112143e+17, 1.282162199212142e+17, 1.282162199312143e+17, 1.282162199412142e+17, 1.282162199512143e+17, 1.282162199612142e+17, 1.282162199712143e+17, 1.282162199812142e+17, 1.282162199912142e+17, 1.282162200012142e+17, 1.282162200112142e+17, 1.282162200212143e+17, 1.282162200312142e+17, 1.282162200412142e+17, 1.282162200512142e+17, 1.282162200612143e+17, 1.282162200712142e+17, 1.282162200812143e+17, 1.282162200912142e+17, 1.282162201012143e+17, 1.282162201112142e+17, 1.282162201212142e+17, 1.282162201312143e+17, 1.282162201412142e+17, 1.282162201512142e+17, 1.282162201612142e+17, 1.282162201712143e+17, 1.282162201812142e+17, 1.282162201912143e+17, 1.282162202012142e+17, 1.282162202112143e+17, 1.282162202212142e+17, 1.282162202312143e+17, 1.282162202412142e+17, 1.282162202512142e+17, 1.282162202612142e+17, 1.282162202712142e+17, 1.282162202812143e+17, 1.282162202912142e+17, 1.282162203012142e+17, 1.282162203112142e+17, 1.282162203212143e+17, 1.282162203312142e+17, 1.282162203412143e+17, 1.282162203512142e+17, 1.282162203612143e+17, 1.282162203712142e+17, 1.282162203812142e+17, 1.282162203912143e+17, 1.282162204012142e+17, 1.282162204112142e+17, 1.282162204212142e+17, 1.282162204312143e+17, 1.282162204412142e+17, 1.282162204512143e+17, 1.282162204612142e+17, 1.282162204712143e+17, 1.282162204812142e+17, 1.282162204912142e+17, 1.282162205012143e+17, 1.282162205112142e+17, 1.282162205212142e+17, 1.282162205312142e+17, 1.282162205412143e+17, 1.282162205512142e+17, 1.282162205612142e+17, 1.282162205712142e+17, 1.282162205812143e+17, 1.282162205912142e+17, 1.282162206012143e+17, 1.282162206112142e+17, 1.282162206212142e+17, 1.282162206312142e+17, 1.282162206412142e+17, 1.282162206512143e+17, 1.282162206612142e+17, 1.282162206712142e+17, 1.282162206812142e+17, 1.282162206912143e+17, 1.282162207012142e+17, 1.282162207112143e+17, 1.282162207212142e+17, 1.282162207312143e+17, 1.282162207412142e+17, 1.282162207512142e+17, 1.282162207612143e+17, 1.282162207712142e+17, 1.282162207812142e+17, 1.282162207912142e+17, 1.282162208012143e+17, 1.282162208112142e+17, 1.282162208212143e+17, 1.282162208312142e+17, 1.282162208412143e+17, 1.282162208512142e+17, 1.282162208612143e+17, 1.282162208712142e+17, 1.282162208812142e+17, 1.282162208912142e+17, 1.282162209012142e+17, 1.282162209112143e+17, 1.282162209212142e+17, 1.282162209312142e+17, 1.282162209412142e+17, 1.282162209512143e+17, 1.282162209612142e+17, 1.282162209712143e+17, 1.282162209812142e+17, 1.282162209912143e+17, 1.282162210012142e+17, 1.282162210112142e+17, 1.282162210212143e+17, 1.282162210312142e+17, 1.282162210412142e+17, 1.282162210512142e+17, 1.282162210612143e+17, 1.282162210712142e+17, 1.282162210812143e+17, 1.282162210912142e+17, 1.282162211012143e+17, 1.282162211112142e+17, 1.282162211212143e+17, 1.282162211312142e+17, 1.282162211412142e+17, 1.282162211512142e+17, 1.282162211612142e+17, 1.282162211712143e+17, 1.282162211812142e+17, 1.282162211912142e+17, 1.282162212012142e+17, 1.282162212112143e+17, 1.282162212212142e+17, 1.282162212312143e+17, 1.282162212412142e+17, 1.282162212512143e+17, 1.282162212612142e+17, 1.282162212712142e+17, 1.282162212812143e+17, 1.282162212912142e+17, 1.282162213012142e+17, 1.282162213112142e+17, 1.282162213212143e+17, 1.282162213312142e+17, 1.282162213412143e+17, 1.282162213512142e+17, 1.282162213612143e+17, 1.282162213712142e+17, 1.282162213812143e+17, 1.282162213912143e+17, 1.282162214012142e+17, 1.282162214112142e+17, 1.282162214212142e+17, 1.282162214312143e+17, 1.282162214412142e+17, 1.282162214512142e+17, 1.282162214612142e+17, 1.282162214712143e+17, 1.282162214812142e+17, 1.282162214912143e+17, 1.282162215012142e+17, 1.282162215112142e+17, 1.282162215212142e+17, 1.282162215312142e+17, 1.282162215412143e+17, 1.282162215512142e+17, 1.282162215612142e+17, 1.282162215712142e+17, 1.282162215812143e+17, 1.282162215912142e+17, 1.282162216012143e+17, 1.282162216112142e+17, 1.282162216212143e+17, 1.282162216312142e+17, 1.282162216412142e+17, 1.282162216512143e+17, 1.282162216612142e+17, 1.282162216712142e+17, 1.282162216812142e+17, 1.282162216912143e+17, 1.282162217012142e+17, 1.282162217112143e+17, 1.282162217212142e+17, 1.282162217312143e+17, 1.282162217412142e+17, 1.282162217512143e+17, 1.282162217612142e+17, 1.282162217712142e+17, 1.282162217812142e+17, 1.282162217912142e+17, 1.282162218012143e+17, 1.282162218112142e+17, 1.282162218212142e+17, 1.282162218312142e+17, 1.282162218412143e+17, 1.282162218512142e+17, 1.282162218612143e+17, 1.282162218712142e+17, 1.282162218812143e+17, 1.282162218912142e+17, 1.282162219012142e+17, 1.282162219112143e+17, 1.282162219212142e+17, 1.282162219312142e+17, 1.282162219412142e+17, 1.282162219512143e+17, 1.282162219612142e+17, 1.282162219712143e+17, 1.282162219812142e+17, 1.282162219912143e+17, 1.282162220012142e+17, 1.282162220112143e+17, 1.282162220212142e+17, 1.282162220312142e+17, 1.282162220412142e+17, 1.282162220512142e+17, 1.282162220612143e+17, 1.282162220712142e+17, 1.282162220812142e+17, 1.282162220912142e+17, 1.282162221012143e+17, 1.282162221112142e+17, 1.282162221212143e+17, 1.282162221312142e+17, 1.282162221412143e+17, 1.282162221512142e+17, 1.282162221612142e+17, 1.282162221712143e+17, 1.282162221812142e+17, 1.282162221912142e+17, 1.282162222012142e+17, 1.282162222112143e+17, 1.282162222212142e+17, 1.282162222312143e+17, 1.282162222412142e+17, 1.282162222512143e+17, 1.282162222612142e+17, 1.282162222712143e+17, 1.282162222812142e+17, 1.282162222912142e+17, 1.282162223012142e+17, 1.282162223112142e+17, 1.282162223212143e+17, 1.282162223312142e+17, 1.282162223412142e+17, 1.282162223512142e+17, 1.282162223612143e+17, 1.282162223712142e+17, 1.282162223812143e+17, 1.282162223912142e+17, 1.282162224012142e+17, 1.282162224112142e+17, 1.282162224212142e+17, 1.282162224312143e+17, 1.282162224412142e+17, 1.282162224512142e+17, 1.282162224612142e+17, 1.282162224712143e+17, 1.282162224812142e+17, 1.282162224912143e+17, 1.282162225012142e+17, 1.282162225112143e+17, 1.282162225212142e+17, 1.282162225312142e+17, 1.282162225412143e+17, 1.282162225512142e+17, 1.282162225612142e+17, 1.282162225712142e+17, 1.282162225812143e+17, 1.282162225912142e+17, 1.282162226012143e+17, 1.282162226112142e+17, 1.282162226212143e+17, 1.282162226312142e+17, 1.282162226412143e+17, 1.282162226512142e+17, 1.282162226612142e+17, 1.282162226712142e+17, 1.282162226812142e+17, 1.282162226912143e+17, 1.282162227012142e+17, 1.282162227112142e+17, 1.282162227212142e+17, 1.282162227312143e+17, 1.282162227412142e+17, 1.282162227512143e+17, 1.282162227612142e+17, 1.282162227712143e+17, 1.282162227812142e+17, 1.282162227912142e+17, 1.282162228012143e+17, 1.282162228112142e+17, 1.282162228212142e+17, 1.282162228312142e+17, 1.282162228412143e+17, 1.282162228512142e+17, 1.282162228612143e+17, 1.282162228712142e+17, 1.282162228812143e+17, 1.282162228912142e+17, 1.282162229012143e+17, 1.282162229112142e+17, 1.282162229212142e+17, 1.282162229312142e+17, 1.282162229412142e+17, 1.282162229512143e+17, 1.282162229612142e+17, 1.282162229712142e+17, 1.282162229812142e+17, 1.282162229912143e+17, 1.282162230012142e+17, 1.282162230112143e+17, 1.282162230212142e+17, 1.282162230312143e+17, 1.282162230412142e+17, 1.282162230512142e+17, 1.282162230612143e+17, 1.282162230712142e+17, 1.282162230812142e+17, 1.282162230912142e+17, 1.282162231012143e+17, 1.282162231112142e+17, 1.282162231212143e+17, 1.282162231312142e+17, 1.282162231412143e+17, 1.282162231512142e+17, 1.282162231612143e+17, 1.282162231712142e+17, 1.282162231812142e+17, 1.282162231912142e+17, 1.282162232012142e+17, 1.282162232112143e+17, 1.282162232212142e+17, 1.282162232312142e+17, 1.282162232412142e+17, 1.282162232512143e+17, 1.282162232612142e+17, 1.282162232712143e+17, 1.282162232812142e+17, 1.282162232912143e+17, 1.282162233012142e+17, 1.282162233112142e+17, 1.282162233212143e+17, 1.282162233312142e+17, 1.282162233412142e+17, 1.282162233512142e+17, 1.282162233612143e+17, 1.282162233712142e+17, 1.282162233812143e+17, 1.282162233912142e+17, 1.282162234012143e+17, 1.282162234112142e+17, 1.282162234212142e+17, 1.282162234312143e+17, 1.282162234412142e+17, 1.282162234512142e+17, 1.282162234612142e+17, 1.282162234712143e+17, 1.282162234812142e+17, 1.282162234912143e+17, 1.282162235012142e+17, 1.282162235112143e+17, 1.282162235212142e+17, 1.282162235312143e+17, 1.282162235412142e+17, 1.282162235512142e+17, 1.282162235612142e+17, 1.282162235712142e+17, 1.282162235812143e+17, 1.282162235912142e+17, 1.282162236012142e+17, 1.282162236112142e+17, 1.282162236212143e+17, 1.282162236312142e+17, 1.282162236412143e+17, 1.282162236512142e+17, 1.282162236612143e+17, 1.282162236712142e+17, 1.282162236812142e+17, 1.282162236912143e+17, 1.282162237012142e+17, 1.282162237112142e+17, 1.282162237212142e+17, 1.282162237312143e+17, 1.282162237412142e+17, 1.282162237512143e+17, 1.282162237612142e+17, 1.282162237712143e+17, 1.282162237812142e+17, 1.282162237912143e+17, 1.282162238012142e+17, 1.282162238112142e+17, 1.282162238212142e+17, 1.282162238312142e+17, 1.282162238412143e+17, 1.282162238512142e+17, 1.282162238612142e+17, 1.282162238712142e+17, 1.282162238812143e+17, 1.282162238912142e+17, 1.282162239012143e+17, 1.282162239112142e+17, 1.282162239212143e+17, 1.282162239312142e+17, 1.282162239412142e+17, 1.282162239512143e+17, 1.282162239612142e+17, 1.282162239712142e+17, 1.282162239812142e+17, 1.282162239912143e+17, 1.282162240012142e+17, 1.282162240112143e+17, 1.282162240212142e+17, 1.282162240312143e+17, 1.282162240412142e+17, 1.282162240512143e+17, 1.282162240612142e+17, 1.282162240712142e+17, 1.282162240812142e+17, 1.282162240912142e+17, 1.282162241012143e+17, 1.282162241112142e+17, 1.282162241212142e+17, 1.282162241312142e+17, 1.282162241412143e+17, 1.282162241512142e+17, 1.282162241612143e+17, 1.282162241712142e+17, 1.282162241812143e+17, 1.282162241912142e+17, 1.282162242012142e+17, 1.282162242112143e+17, 1.282162242212142e+17, 1.282162242312142e+17, 1.282162242412142e+17, 1.282162242512143e+17, 1.282162242612142e+17, 1.282162242712143e+17, 1.282162242812142e+17, 1.282162242912143e+17, 1.282162243012142e+17, 1.282162243112142e+17, 1.282162243212143e+17, 1.282162243312142e+17, 1.282162243412142e+17, 1.282162243512142e+17, 1.282162243612143e+17, 1.282162243712142e+17, 1.282162243812142e+17, 1.282162243912142e+17, 1.282162244012143e+17, 1.282162244112142e+17, 1.282162244212143e+17, 1.282162244312142e+17, 1.282162244412142e+17, 1.282162244512142e+17, 1.282162244612142e+17, 1.282162244712143e+17, 1.282162244812142e+17, 1.282162244912142e+17, 1.282162245012142e+17, 1.282162245112143e+17, 1.282162245212142e+17, 1.282162245312143e+17, 1.282162245412142e+17, 1.282162245512143e+17, 1.282162245612142e+17, 1.282162245712142e+17, 1.282162245812143e+17, 1.282162245912142e+17, 1.282162246012142e+17, 1.282162246112142e+17, 1.282162246212143e+17, 1.282162246312142e+17, 1.282162246412143e+17, 1.282162246512142e+17, 1.282162246612143e+17, 1.282162246712142e+17, 1.282162246812143e+17, 1.282162246912142e+17, 1.282162247012142e+17, 1.282162247112142e+17, 1.282162247212142e+17, 1.282162247312143e+17, 1.282162247412142e+17, 1.282162247512142e+17, 1.282162247612142e+17, 1.282162247712143e+17, 1.282162247812142e+17, 1.282162247912143e+17, 1.282162248012142e+17, 1.282162248112143e+17, 1.282162248212142e+17, 1.282162248312142e+17, 1.282162248412143e+17, 1.282162248512142e+17, 1.282162248612142e+17, 1.282162248712142e+17, 1.282162248812143e+17, 1.282162248912142e+17, 1.282162249012143e+17, 1.282162249112142e+17, 1.282162249212143e+17, 1.282162249312142e+17, 1.282162249412143e+17, 1.282162249512142e+17, 1.282162249612142e+17, 1.282162249712142e+17, 1.282162249812142e+17, 1.282162249912143e+17, 1.282162250012142e+17, 1.282162250112142e+17, 1.282162250212142e+17, 1.282162250312143e+17, 1.282162250412142e+17, 1.282162250512143e+17, 1.282162250612142e+17, 1.282162250712143e+17, 1.282162250812142e+17, 1.282162250912142e+17, 1.282162251012143e+17, 1.282162251112142e+17, 1.282162251212142e+17, 1.282162251312142e+17, 1.282162251412143e+17, 1.282162251512142e+17, 1.282162251612143e+17, 1.282162251712142e+17, 1.282162251812143e+17, 1.282162251912142e+17, 1.282162252012143e+17, 1.282162252112143e+17, 1.282162252212142e+17, 1.282162252312142e+17, 1.282162252412142e+17, 1.282162252512143e+17, 1.282162252612142e+17, 1.282162252712142e+17, 1.282162252812142e+17, 1.282162252912143e+17, 1.282162253012142e+17, 1.282162253112143e+17, 1.282162253212142e+17, 1.282162253312142e+17, 1.282162253412142e+17, 1.282162253512142e+17, 1.282162253612143e+17, 1.282162253712142e+17, 1.282162253812142e+17, 1.282162253912142e+17, 1.282162254012143e+17, 1.282162254112142e+17, 1.282162254212143e+17, 1.282162254312142e+17, 1.282162254412143e+17, 1.282162254512142e+17, 1.282162254612142e+17, 1.282162254712143e+17, 1.282162254812142e+17, 1.282162254912142e+17, 1.282162255012142e+17, 1.282162255112143e+17, 1.282162255212142e+17, 1.282162255312143e+17, 1.282162255412142e+17, 1.282162255512143e+17, 1.282162255612142e+17, 1.282162255712143e+17, 1.282162255812142e+17, 1.282162255912142e+17, 1.282162256012142e+17, 1.282162256112142e+17, 1.282162256212143e+17, 1.282162256312142e+17, 1.282162256412142e+17, 1.282162256512142e+17, 1.282162256612143e+17, 1.282162256712142e+17, 1.282162256812143e+17, 1.282162256912142e+17, 1.282162257012143e+17, 1.282162257112142e+17, 1.282162257212142e+17, 1.282162257312143e+17, 1.282162257412142e+17, 1.282162257512142e+17, 1.282162257612142e+17, 1.282162257712143e+17, 1.282162257812142e+17, 1.282162257912143e+17, 1.282162258012142e+17, 1.282162258112143e+17, 1.282162258212142e+17, 1.282162258312143e+17, 1.282162258412142e+17, 1.282162258512142e+17, 1.282162258612142e+17, 1.282162258712142e+17, 1.282162258812143e+17, 1.282162258912142e+17, 1.282162259012142e+17, 1.282162259112142e+17, 1.282162259212143e+17, 1.282162259312142e+17, 1.282162259412143e+17, 1.282162259512142e+17, 1.282162259612143e+17, 1.282162259712142e+17, 1.282162259812142e+17, 1.282162259912143e+17, 1.282162260012142e+17, 1.282162260112142e+17, 1.282162260212142e+17, 1.282162260312143e+17, 1.282162260412142e+17, 1.282162260512143e+17, 1.282162260612142e+17, 1.282162260712143e+17, 1.282162260812142e+17, 1.282162260912143e+17, 1.282162261012142e+17, 1.282162261112142e+17, 1.282162261212142e+17, 1.282162261312142e+17, 1.282162261412143e+17, 1.282162261512142e+17, 1.282162261612142e+17, 1.282162261712142e+17, 1.282162261812143e+17, 1.282162261912142e+17, 1.282162262012143e+17, 1.282162262112142e+17, 1.282162262212143e+17, 1.282162262312142e+17, 1.282162262412142e+17, 1.282162262512143e+17, 1.282162262612142e+17, 1.282162262712142e+17, 1.282162262812142e+17, 1.282162262912143e+17, 1.282162263012142e+17, 1.282162263112143e+17, 1.282162263212142e+17, 1.282162263312143e+17, 1.282162263412142e+17, 1.282162263512142e+17, 1.282162263612143e+17, 1.282162263712142e+17, 1.282162263812142e+17, 1.282162263912142e+17, 1.282162264012143e+17, 1.282162264112142e+17, 1.282162264212143e+17, 1.282162264312142e+17, 1.282162264412143e+17, 1.282162264512142e+17, 1.282162264612143e+17, 1.282162264712142e+17, 1.282162264812142e+17},
			             {1.282161925512142e+17, 1.282161925612143e+17, 1.282161925712142e+17, 1.282161925812143e+17, 1.282161925912142e+17, 1.282161926012142e+17, 1.282161926112143e+17, 1.282161926212142e+17, 1.282161926312142e+17, 1.282161926412142e+17, 1.282161926512143e+17, 1.282161926612142e+17, 1.282161926712143e+17, 1.282161926812142e+17, 1.282161926912143e+17, 1.282161927012142e+17, 1.282161927112143e+17, 1.282161927212142e+17, 1.282161927312142e+17, 1.282161927412142e+17, 1.282161927512142e+17, 1.282161927612143e+17, 1.282161927712142e+17, 1.282161927812142e+17, 1.282161927912142e+17, 1.282161928012143e+17, 1.282161928112142e+17, 1.282161928212143e+17, 1.282161928312142e+17, 1.282161928412143e+17, 1.282161928512142e+17, 1.282161928612142e+17, 1.282161928712143e+17, 1.282161928812142e+17, 1.282161928912142e+17, 1.282161929012142e+17, 1.282161929112143e+17, 1.282161929212142e+17, 1.282161929312143e+17, 1.282161929412142e+17, 1.282161929512143e+17, 1.282161929612142e+17, 1.282161929712143e+17, 1.282161929812142e+17, 1.282161929912142e+17, 1.282161930012142e+17, 1.282161930112142e+17, 1.282161930212143e+17, 1.282161930312142e+17, 1.282161930412142e+17, 1.282161930512142e+17, 1.282161930612143e+17, 1.282161930712142e+17, 1.282161930812143e+17, 1.282161930912142e+17, 1.282161931012143e+17, 1.282161931112142e+17, 1.282161931212142e+17, 1.282161931312143e+17, 1.282161931412142e+17, 1.282161931512142e+17, 1.282161931612142e+17, 1.282161931712143e+17, 1.282161931812142e+17, 1.282161931912143e+17, 1.282161932012142e+17, 1.282161932112143e+17, 1.282161932212142e+17, 1.282161932312143e+17, 1.282161932412142e+17, 1.282161932512142e+17, 1.282161932612142e+17, 1.282161932712142e+17, 1.282161932812143e+17, 1.282161932912142e+17, 1.282161933012142e+17, 1.282161933112142e+17, 1.282161933212143e+17, 1.282161933312142e+17, 1.282161933412143e+17, 1.282161933512142e+17, 1.282161933612143e+17, 1.282161933712142e+17, 1.282161933812142e+17, 1.282161933912143e+17, 1.282161934012142e+17, 1.282161934112142e+17, 1.282161934212142e+17, 1.282161934312143e+17, 1.282161934412142e+17, 1.282161934512143e+17, 1.282161934612142e+17, 1.282161934712143e+17, 1.282161934812142e+17, 1.282161934912142e+17, 1.282161935012143e+17, 1.282161935112142e+17, 1.282161935212142e+17, 1.282161935312142e+17, 1.282161935412143e+17, 1.282161935512142e+17, 1.282161935612142e+17, 1.282161935712142e+17, 1.282161935812143e+17, 1.282161935912142e+17, 1.282161936012143e+17, 1.282161936112142e+17, 1.282161936212142e+17, 1.282161936312142e+17, 1.282161936412142e+17, 1.282161936512143e+17, 1.282161936612142e+17, 1.282161936712142e+17, 1.282161936812142e+17, 1.282161936912143e+17, 1.282161937012142e+17, 1.282161937112143e+17, 1.282161937212142e+17, 1.282161937312143e+17, 1.282161937412142e+17, 1.282161937512142e+17, 1.282161937612143e+17, 1.282161937712142e+17, 1.282161937812142e+17, 1.282161937912142e+17, 1.282161938012143e+17, 1.282161938112142e+17, 1.282161938212143e+17, 1.282161938312142e+17, 1.282161938412143e+17, 1.282161938512142e+17, 1.282161938612143e+17, 1.282161938712142e+17, 1.282161938812142e+17, 1.282161938912142e+17, 1.282161939012142e+17, 1.282161939112143e+17, 1.282161939212142e+17, 1.282161939312142e+17, 1.282161939412142e+17, 1.282161939512143e+17, 1.282161939612142e+17, 1.282161939712143e+17, 1.282161939812142e+17, 1.282161939912143e+17, 1.282161940012142e+17, 1.282161940112142e+17, 1.282161940212143e+17, 1.282161940312142e+17, 1.282161940412142e+17, 1.282161940512142e+17, 1.282161940612143e+17, 1.282161940712142e+17, 1.282161940812143e+17, 1.282161940912142e+17, 1.282161941012143e+17, 1.282161941112142e+17, 1.282161941212143e+17, 1.282161941312142e+17, 1.282161941412142e+17, 1.282161941512142e+17, 1.282161941612142e+17, 1.282161941712143e+17, 1.282161941812142e+17, 1.282161941912142e+17, 1.282161942012142e+17, 1.282161942112143e+17, 1.282161942212142e+17, 1.282161942312143e+17, 1.282161942412142e+17, 1.282161942512143e+17, 1.282161942612142e+17, 1.282161942712142e+17, 1.282161942812143e+17, 1.282161942912142e+17, 1.282161943012142e+17, 1.282161943112142e+17, 1.282161943212143e+17, 1.282161943312142e+17, 1.282161943412143e+17, 1.282161943512142e+17, 1.282161943612143e+17, 1.282161943712142e+17, 1.282161943812143e+17, 1.282161943912143e+17, 1.282161944012142e+17, 1.282161944112142e+17, 1.282161944212142e+17, 1.282161944312143e+17, 1.282161944412142e+17, 1.282161944512142e+17, 1.282161944612142e+17, 1.282161944712143e+17, 1.282161944812142e+17, 1.282161944912143e+17, 1.282161945012142e+17, 1.282161945112142e+17, 1.282161945212142e+17, 1.282161945312142e+17, 1.282161945412143e+17, 1.282161945512142e+17, 1.282161945612142e+17, 1.282161945712142e+17, 1.282161945812143e+17, 1.282161945912142e+17, 1.282161946012143e+17, 1.282161946112142e+17, 1.282161946212143e+17, 1.282161946312142e+17, 1.282161946412142e+17, 1.282161946512143e+17, 1.282161946612142e+17, 1.282161946712142e+17, 1.282161946812142e+17, 1.282161946912143e+17, 1.282161947012142e+17, 1.282161947112143e+17, 1.282161947212142e+17, 1.282161947312143e+17, 1.282161947412142e+17, 1.282161947512143e+17, 1.282161947612142e+17, 1.282161947712142e+17, 1.282161947812142e+17, 1.282161947912142e+17, 1.282161948012143e+17, 1.282161948112142e+17, 1.282161948212142e+17, 1.282161948312142e+17, 1.282161948412143e+17, 1.282161948512142e+17, 1.282161948612143e+17, 1.282161948712142e+17, 1.282161948812143e+17, 1.282161948912142e+17, 1.282161949012142e+17, 1.282161949112143e+17, 1.282161949212142e+17, 1.282161949312142e+17, 1.282161949412142e+17, 1.282161949512143e+17, 1.282161949612142e+17, 1.282161949712143e+17, 1.282161949812142e+17, 1.282161949912143e+17, 1.282161950012142e+17, 1.282161950112143e+17, 1.282161950212142e+17, 1.282161950312142e+17, 1.282161950412142e+17, 1.282161950512142e+17, 1.282161950612143e+17, 1.282161950712142e+17, 1.282161950812142e+17, 1.282161950912142e+17, 1.282161951012143e+17, 1.282161951112142e+17, 1.282161951212143e+17, 1.282161951312142e+17, 1.282161951412143e+17, 1.282161951512142e+17, 1.282161951612142e+17, 1.282161951712143e+17, 1.282161951812142e+17, 1.282161951912142e+17, 1.282161952012142e+17, 1.282161952112143e+17, 1.282161952212142e+17, 1.282161952312143e+17, 1.282161952412142e+17, 1.282161952512143e+17, 1.282161952612142e+17, 1.282161952712143e+17, 1.282161952812142e+17, 1.282161952912142e+17, 1.282161953012142e+17, 1.282161953112142e+17, 1.282161953212143e+17, 1.282161953312142e+17, 1.282161953412142e+17, 1.282161953512142e+17, 1.282161953612143e+17, 1.282161953712142e+17, 1.282161953812143e+17, 1.282161953912142e+17, 1.282161954012142e+17, 1.282161954112142e+17, 1.282161954212142e+17, 1.282161954312143e+17, 1.282161954412142e+17, 1.282161954512142e+17, 1.282161954612142e+17, 1.282161954712143e+17, 1.282161954812142e+17, 1.282161954912143e+17, 1.282161955012142e+17, 1.282161955112143e+17, 1.282161955212142e+17, 1.282161955312142e+17, 1.282161955412143e+17, 1.282161955512142e+17, 1.282161955612142e+17, 1.282161955712142e+17, 1.282161955812143e+17, 1.282161955912142e+17, 1.282161956012143e+17, 1.282161956112142e+17, 1.282161956212143e+17, 1.282161956312142e+17, 1.282161956412143e+17, 1.282161956512142e+17, 1.282161956612142e+17, 1.282161956712142e+17, 1.282161956812142e+17, 1.282161956912143e+17, 1.282161957012142e+17, 1.282161957112142e+17, 1.282161957212142e+17, 1.282161957312143e+17, 1.282161957412142e+17, 1.282161957512143e+17, 1.282161957612142e+17, 1.282161957712143e+17, 1.282161957812142e+17, 1.282161957912142e+17, 1.282161958012143e+17, 1.282161958112142e+17, 1.282161958212142e+17, 1.282161958312142e+17, 1.282161958412143e+17, 1.282161958512142e+17, 1.282161958612143e+17, 1.282161958913705e+17, 1.282161959012143e+17, 1.282161959112142e+17, 1.282161959212142e+17, 1.282161959312142e+17, 1.282161959512143e+17, 1.282161959612142e+17, 1.282161959712142e+17, 1.282161959812142e+17, 1.282161959912143e+17, 1.282161960012142e+17, 1.282161960112143e+17, 1.282161960212142e+17, 1.282161960312143e+17, 1.282161960412142e+17, 1.282161960512142e+17, 1.282161960612143e+17, 1.282161960712142e+17, 1.282161960812142e+17, 1.282161960912142e+17, 1.282161961012143e+17, 1.282161961112142e+17, 1.282161961212143e+17, 1.282161961312142e+17, 1.282161961412143e+17, 1.282161961512142e+17, 1.282161961612143e+17, 1.282161961712142e+17, 1.282161961812142e+17, 1.282161961912142e+17, 1.282161962012142e+17, 1.282161962112143e+17, 1.282161962212142e+17, 1.282161962312142e+17, 1.282161962412142e+17, 1.282161962512143e+17, 1.282161962612142e+17, 1.282161962712143e+17, 1.282161962812142e+17, 1.282161962912143e+17, 1.282161963012142e+17, 1.282161963112142e+17, 1.282161963212143e+17, 1.282161963312142e+17, 1.282161963412142e+17, 1.282161963512142e+17, 1.282161963612143e+17, 1.282161963712142e+17, 1.282161963812143e+17, 1.282161963912142e+17, 1.282161964012143e+17, 1.282161964112142e+17, 1.282161964212142e+17, 1.282161964312143e+17, 1.282161964412142e+17, 1.282161964512142e+17, 1.282161964612142e+17, 1.282161964712143e+17, 1.282161964812142e+17, 1.282161964912143e+17, 1.282161965012142e+17, 1.282161965112143e+17, 1.282161965212142e+17, 1.282161965312143e+17, 1.282161965412142e+17, 1.282161965512142e+17, 1.282161965612142e+17, 1.282161965712142e+17, 1.282161965812143e+17, 1.282161965912142e+17, 1.282161966012142e+17, 1.282161966112142e+17, 1.282161966212143e+17, 1.282161966312142e+17, 1.282161966412143e+17, 1.282161966512142e+17, 1.282161966612143e+17, 1.282161966712142e+17, 1.282161966812142e+17, 1.282161966912143e+17, 1.282161967012142e+17, 1.282161967112142e+17, 1.282161967212142e+17, 1.282161967312143e+17, 1.282161967412142e+17, 1.282161967512143e+17, 1.282161967612142e+17, 1.282161967712143e+17, 1.282161967812142e+17, 1.282161967912143e+17, 1.282161968012142e+17, 1.282161968112142e+17, 1.282161968212142e+17, 1.282161968312142e+17, 1.282161968412143e+17, 1.282161968512142e+17, 1.282161968612142e+17, 1.282161968712142e+17, 1.282161968812143e+17, 1.282161968912142e+17, 1.282161969012143e+17, 1.282161969112142e+17, 1.282161969212143e+17, 1.282161969312142e+17, 1.282161969412142e+17, 1.282161969512143e+17, 1.282161969612142e+17, 1.282161969712142e+17, 1.282161969812142e+17, 1.282161969912143e+17, 1.282161970012142e+17, 1.282161970112143e+17, 1.282161970212142e+17, 1.282161970312143e+17, 1.282161970412142e+17, 1.282161970512143e+17, 1.282161970612142e+17, 1.282161970712142e+17, 1.282161970812142e+17, 1.282161970912142e+17, 1.282161971012143e+17, 1.282161971112142e+17, 1.282161971212142e+17, 1.282161971312142e+17, 1.282161971412143e+17, 1.282161971512142e+17, 1.282161971612143e+17, 1.282161971712142e+17, 1.282161971812143e+17, 1.282161971912142e+17, 1.282161972012142e+17, 1.282161972112143e+17, 1.282161972212142e+17, 1.282161972312142e+17, 1.282161972412142e+17, 1.282161972512143e+17, 1.282161972612142e+17, 1.282161972712143e+17, 1.282161972812142e+17, 1.282161972912143e+17, 1.282161973012142e+17, 1.282161973112142e+17, 1.282161973212143e+17, 1.282161973312142e+17, 1.282161973412142e+17, 1.282161973512142e+17, 1.282161973612143e+17, 1.282161973712142e+17, 1.282161973812142e+17, 1.282161973912142e+17, 1.282161974012143e+17, 1.282161974112142e+17, 1.282161974212143e+17, 1.282161974312142e+17, 1.282161974412142e+17, 1.282161974512142e+17, 1.282161974612142e+17, 1.282161974712143e+17, 1.282161974812142e+17, 1.282161974912142e+17, 1.282161975012142e+17, 1.282161975112143e+17, 1.282161975212142e+17, 1.282161975312143e+17, 1.282161975412142e+17, 1.282161975512143e+17, 1.282161975612142e+17, 1.282161975712142e+17, 1.282161975812143e+17, 1.282161975912142e+17, 1.282161976012142e+17, 1.282161976112142e+17, 1.282161976212143e+17, 1.282161976312142e+17, 1.282161976412143e+17, 1.282161976512142e+17, 1.282161976612143e+17, 1.282161976712142e+17, 1.282161976812143e+17, 1.282161976912142e+17, 1.282161977012142e+17, 1.282161977112142e+17, 1.282161977212142e+17, 1.282161977312143e+17, 1.282161977412142e+17, 1.282161977512142e+17, 1.282161977612142e+17, 1.282161977712143e+17, 1.282161977812142e+17, 1.282161977912143e+17, 1.282161978012142e+17, 1.282161978112143e+17, 1.282161978212142e+17, 1.282161978312142e+17, 1.282161978412143e+17, 1.282161978512142e+17, 1.282161978612142e+17, 1.282161978712142e+17, 1.282161978812143e+17, 1.282161978912142e+17, 1.282161979012143e+17, 1.282161979112142e+17, 1.282161979212143e+17, 1.282161979312142e+17, 1.282161979412143e+17, 1.282161979512142e+17, 1.282161979612142e+17, 1.282161979712142e+17, 1.282161979812142e+17, 1.282161979912143e+17, 1.282161980012142e+17, 1.282161980112142e+17, 1.282161980212142e+17, 1.282161980312143e+17, 1.282161980412142e+17, 1.282161980512143e+17, 1.282161980612142e+17, 1.282161980712143e+17, 1.282161980812142e+17, 1.282161980912142e+17, 1.282161981012143e+17, 1.282161981112142e+17, 1.282161981212142e+17, 1.282161981312142e+17, 1.282161981412143e+17, 1.282161981512142e+17, 1.282161981612143e+17, 1.282161981712142e+17, 1.282161981812143e+17, 1.282161981912142e+17, 1.282161982012143e+17, 1.282161982112143e+17, 1.282161982212142e+17, 1.282161982312142e+17, 1.282161982412142e+17, 1.282161982512143e+17, 1.282161982612142e+17, 1.282161982712142e+17, 1.282161982812142e+17, 1.282161982912143e+17, 1.282161983012142e+17, 1.282161983112143e+17, 1.282161983212142e+17, 1.282161983312142e+17, 1.282161983412142e+17, 1.282161983512142e+17, 1.282161983612143e+17, 1.282161983712142e+17, 1.282161983812142e+17, 1.282161983912142e+17, 1.282161984012143e+17, 1.282161984112142e+17, 1.282161984212143e+17, 1.282161984312142e+17, 1.282161984412143e+17, 1.282161984512142e+17, 1.282161984612142e+17, 1.282161984712143e+17, 1.282161984812142e+17, 1.282161984912142e+17, 1.282161985012142e+17, 1.282161985112143e+17, 1.282161985212142e+17, 1.282161985312143e+17, 1.282161985412142e+17, 1.282161985512143e+17, 1.282161985612142e+17, 1.282161985712143e+17, 1.282161985812142e+17, 1.282161985912142e+17, 1.282161986012142e+17, 1.282161986112142e+17, 1.282161986212143e+17, 1.282161986312142e+17, 1.282161986412142e+17, 1.282161986512142e+17, 1.282161986612143e+17, 1.282161986712142e+17, 1.282161986812143e+17, 1.282161986912142e+17, 1.282161987012143e+17, 1.282161987112142e+17, 1.282161987212142e+17, 1.282161987312143e+17, 1.282161987412142e+17, 1.282161987512142e+17, 1.282161987612142e+17, 1.282161987712143e+17, 1.282161987812142e+17, 1.282161987912143e+17, 1.282161988012142e+17, 1.282161988112143e+17, 1.282161988212142e+17, 1.282161988312143e+17, 1.282161988412142e+17, 1.282161988512142e+17, 1.282161988612142e+17, 1.282161988712142e+17, 1.282161988812143e+17, 1.282161988912142e+17, 1.282161989012142e+17, 1.282161989112142e+17, 1.282161989212143e+17, 1.282161989312142e+17, 1.282161989412143e+17, 1.282161989512142e+17, 1.282161989612143e+17, 1.282161989712142e+17, 1.282161989812142e+17, 1.282161989912143e+17, 1.282161990012142e+17, 1.282161990112142e+17, 1.282161990212142e+17, 1.282161990312143e+17, 1.282161990412142e+17, 1.282161990512143e+17, 1.282161990612142e+17, 1.282161990712143e+17, 1.282161990812142e+17, 1.282161990912143e+17, 1.282161991012142e+17, 1.282161991112142e+17, 1.282161991212142e+17, 1.282161991312142e+17, 1.282161991412143e+17, 1.282161991512142e+17, 1.282161991612142e+17, 1.282161991712142e+17, 1.282161991812143e+17, 1.282161991912142e+17, 1.282161992012143e+17, 1.282161992112142e+17, 1.282161992212143e+17, 1.282161992312142e+17, 1.282161992412142e+17, 1.282161992512143e+17, 1.282161992612142e+17, 1.282161992712142e+17, 1.282161992812142e+17, 1.282161992912143e+17, 1.282161993012142e+17, 1.282161993112143e+17, 1.282161993212142e+17, 1.282161993312143e+17, 1.282161993412142e+17, 1.282161993512142e+17, 1.282161993612143e+17, 1.282161993712142e+17, 1.282161993812142e+17, 1.282161993912142e+17, 1.282161994012143e+17, 1.282161994112142e+17, 1.282161994212143e+17, 1.282161994312142e+17, 1.282161994412143e+17, 1.282161994512142e+17, 1.282161994612143e+17, 1.282161994712142e+17, 1.282161994812142e+17, 1.282161994912142e+17, 1.282161995012142e+17, 1.282161995112143e+17, 1.282161995212142e+17, 1.282161995312142e+17, 1.282161995412142e+17, 1.282161995512143e+17, 1.282161995612142e+17, 1.282161995712143e+17, 1.282161995812142e+17, 1.282161995912143e+17, 1.282161996012142e+17, 1.282161996112142e+17, 1.282161996212143e+17, 1.282161996312142e+17, 1.282161996412142e+17, 1.282161996512142e+17, 1.282161996612143e+17, 1.282161996712142e+17, 1.282161996812143e+17, 1.282161996912142e+17, 1.282161997012143e+17, 1.282161997112142e+17, 1.282161997212143e+17, 1.282161997312142e+17, 1.282161997412142e+17, 1.282161997512142e+17, 1.282161997612142e+17, 1.282161997712143e+17, 1.282161997812142e+17, 1.282161997912142e+17, 1.282161998012142e+17, 1.282161998112143e+17, 1.282161998212142e+17, 1.282161998312143e+17, 1.282161998412142e+17, 1.282161998512143e+17, 1.282161998612142e+17, 1.282161998712142e+17, 1.282161998812143e+17, 1.282161998912142e+17, 1.282161999012142e+17, 1.282161999112142e+17, 1.282161999212143e+17, 1.282161999312142e+17, 1.282161999412143e+17, 1.282161999512142e+17, 1.282161999612143e+17, 1.282161999712142e+17, 1.282161999812143e+17, 1.282161999912142e+17, 1.282162000012142e+17, 1.282162000112142e+17, 1.282162000212142e+17, 1.282162000312143e+17, 1.282162000412142e+17, 1.282162000512142e+17, 1.282162000612142e+17, 1.282162000712143e+17, 1.282162000812142e+17, 1.282162000912143e+17, 1.282162001012142e+17, 1.282162001112143e+17, 1.282162001212142e+17, 1.282162001312142e+17, 1.282162001412143e+17, 1.282162001512142e+17, 1.282162001612142e+17, 1.282162001712142e+17, 1.282162001812143e+17, 1.282162001912142e+17, 1.282162002012143e+17, 1.282162002112142e+17, 1.282162002212143e+17, 1.282162002312142e+17, 1.282162002412142e+17, 1.282162002512143e+17, 1.282162002612142e+17, 1.282162002712142e+17, 1.282162002812142e+17, 1.282162002912143e+17, 1.282162003012142e+17, 1.282162003112142e+17, 1.282162003212142e+17, 1.282162003312143e+17, 1.282162003412142e+17, 1.282162003512143e+17, 1.282162003612142e+17, 1.282162003712142e+17, 1.282162003812142e+17, 1.282162003912142e+17, 1.282162004012143e+17, 1.282162004112142e+17, 1.282162004212142e+17, 1.282162004312142e+17, 1.282162004412143e+17, 1.282162004512142e+17, 1.282162004612143e+17, 1.282162004712142e+17, 1.282162004812143e+17, 1.282162004912142e+17, 1.282162005012142e+17, 1.282162005112143e+17, 1.282162005212142e+17, 1.282162005312142e+17, 1.282162005412142e+17, 1.282162005512143e+17, 1.282162005612142e+17, 1.282162005712143e+17, 1.282162005812142e+17, 1.282162005912143e+17, 1.282162006012142e+17, 1.282162006112143e+17, 1.282162006212142e+17, 1.282162006312142e+17, 1.282162006412142e+17, 1.282162006512142e+17, 1.282162006612143e+17, 1.282162006712142e+17, 1.282162006812142e+17, 1.282162006912142e+17, 1.282162007012143e+17, 1.282162007112142e+17, 1.282162007212143e+17, 1.282162007312142e+17, 1.282162007412143e+17, 1.282162007512142e+17, 1.282162007612142e+17, 1.282162007712143e+17, 1.282162007812142e+17, 1.282162007912142e+17, 1.282162008012142e+17, 1.282162008112143e+17, 1.282162008212142e+17, 1.282162008312143e+17, 1.282162008412142e+17, 1.282162008512143e+17, 1.282162008612142e+17, 1.282162008712143e+17, 1.282162008812142e+17, 1.282162008912142e+17, 1.282162009012142e+17, 1.282162009112142e+17, 1.282162009212143e+17, 1.282162009312142e+17, 1.282162009412142e+17, 1.282162009512142e+17, 1.282162009612143e+17, 1.282162009712142e+17, 1.282162009812143e+17, 1.282162009912142e+17, 1.282162010012143e+17, 1.282162010112142e+17, 1.282162010212142e+17, 1.282162010312143e+17, 1.282162010412142e+17, 1.282162010512142e+17, 1.282162010612142e+17, 1.282162010712143e+17, 1.282162010812142e+17, 1.282162010912143e+17, 1.282162011012142e+17, 1.282162011112143e+17, 1.282162011212142e+17, 1.282162011312143e+17, 1.282162011412143e+17, 1.282162011512142e+17, 1.282162011612142e+17, 1.282162011712142e+17, 1.282162011812143e+17, 1.282162011912142e+17, 1.282162012012142e+17, 1.282162012112142e+17, 1.282162012212143e+17, 1.282162012312142e+17, 1.282162012412143e+17, 1.282162012512142e+17, 1.282162012612142e+17, 1.282162012712142e+17, 1.282162012812142e+17, 1.282162012912143e+17, 1.282162013012142e+17, 1.282162013112142e+17, 1.282162013212142e+17, 1.282162013312143e+17, 1.282162013412142e+17, 1.282162013512143e+17, 1.282162013612142e+17, 1.282162013712143e+17, 1.282162013812142e+17, 1.282162013912142e+17, 1.282162014012143e+17, 1.282162014112142e+17, 1.282162014212142e+17, 1.282162014312142e+17, 1.282162014412143e+17, 1.282162014512142e+17, 1.282162014612143e+17, 1.282162014712142e+17, 1.282162014812143e+17, 1.282162014912142e+17, 1.282162015012143e+17, 1.282162015112142e+17, 1.282162015212142e+17, 1.282162015312142e+17, 1.282162015412142e+17, 1.282162015512143e+17, 1.282162015612142e+17, 1.282162015712142e+17, 1.282162015812142e+17, 1.282162015912143e+17, 1.282162016012142e+17, 1.282162016112143e+17, 1.282162016212142e+17, 1.282162016312143e+17, 1.282162016412142e+17, 1.282162016512142e+17, 1.282162016612143e+17, 1.282162016712142e+17, 1.282162016812142e+17, 1.282162016912142e+17, 1.282162017012143e+17, 1.282162017112142e+17, 1.282162017212143e+17, 1.282162017312142e+17, 1.282162017412143e+17, 1.282162017512142e+17, 1.282162017612143e+17, 1.282162017712142e+17, 1.282162017812142e+17, 1.282162017912142e+17, 1.282162018012142e+17, 1.282162018112143e+17, 1.282162018212142e+17, 1.282162018312142e+17, 1.282162018412142e+17, 1.282162018512143e+17, 1.282162018612142e+17, 1.282162018712143e+17, 1.282162018812142e+17, 1.282162018912143e+17, 1.282162019012142e+17, 1.282162019112142e+17, 1.282162019212143e+17, 1.282162019312142e+17, 1.282162019412142e+17, 1.282162019512142e+17, 1.282162019612143e+17, 1.282162019712142e+17, 1.282162019812143e+17, 1.282162019912142e+17, 1.282162020012143e+17, 1.282162020112142e+17, 1.282162020212143e+17, 1.282162020312142e+17, 1.282162020412142e+17, 1.282162020512142e+17, 1.282162020612142e+17, 1.282162020712143e+17, 1.282162020812142e+17, 1.282162020912142e+17, 1.282162021012142e+17, 1.282162021112143e+17, 1.282162021212142e+17, 1.282162021312143e+17, 1.282162021412142e+17, 1.282162021512142e+17, 1.282162021612142e+17, 1.282162021712142e+17, 1.282162021812143e+17, 1.282162021912142e+17, 1.282162022012142e+17, 1.282162022112142e+17, 1.282162022212143e+17, 1.282162022312142e+17, 1.282162022412143e+17, 1.282162022512142e+17, 1.282162022612143e+17, 1.282162022712142e+17, 1.282162022812142e+17, 1.282162022912143e+17, 1.282162023012142e+17, 1.282162023112142e+17, 1.282162023212142e+17, 1.282162023312143e+17, 1.282162023412142e+17, 1.282162023512143e+17, 1.282162023612142e+17, 1.282162023712143e+17, 1.282162023812142e+17, 1.282162023912143e+17, 1.282162024012142e+17, 1.282162024112142e+17, 1.282162024212142e+17, 1.282162024312142e+17, 1.282162024412143e+17, 1.282162024512142e+17, 1.282162024612142e+17, 1.282162024712142e+17, 1.282162024812143e+17, 1.282162024912142e+17, 1.282162025012143e+17, 1.282162025112142e+17, 1.282162025212143e+17, 1.282162025312142e+17, 1.282162025412142e+17, 1.282162025512143e+17, 1.282162025612142e+17, 1.282162025712142e+17, 1.282162025812142e+17, 1.282162025912143e+17, 1.282162026012142e+17, 1.282162026112143e+17, 1.282162026212142e+17, 1.282162026312143e+17, 1.282162026412142e+17, 1.282162026512143e+17, 1.282162026612142e+17, 1.282162026712142e+17, 1.282162026812142e+17, 1.282162026912142e+17, 1.282162027012143e+17, 1.282162027112142e+17, 1.282162027212142e+17, 1.282162027312142e+17, 1.282162027412143e+17, 1.282162027512142e+17, 1.282162027612143e+17, 1.282162027712142e+17, 1.282162027812143e+17, 1.282162027912142e+17, 1.282162028012142e+17, 1.282162028112143e+17, 1.282162028212142e+17, 1.282162028312142e+17, 1.282162028412142e+17, 1.282162028512143e+17, 1.282162028612142e+17, 1.282162028712143e+17, 1.282162028812142e+17, 1.282162028912143e+17, 1.282162029012142e+17, 1.282162029112143e+17, 1.282162029212142e+17, 1.282162029312142e+17, 1.282162029412142e+17, 1.282162029512142e+17, 1.282162029612143e+17, 1.282162029712142e+17, 1.282162029812142e+17, 1.282162029912142e+17, 1.282162030012143e+17, 1.282162030112142e+17, 1.282162030212143e+17, 1.282162030312142e+17, 1.282162030412143e+17, 1.282162030512142e+17, 1.282162030612142e+17, 1.282162030712143e+17, 1.282162030812142e+17, 1.282162030912142e+17, 1.282162031012142e+17, 1.282162031112143e+17, 1.282162031212142e+17, 1.282162031312143e+17, 1.282162031412142e+17, 1.282162031512143e+17, 1.282162031612142e+17, 1.282162031712142e+17, 1.282162031812143e+17, 1.282162031912142e+17, 1.282162032012142e+17, 1.282162032112142e+17, 1.282162032212143e+17, 1.282162032312142e+17, 1.282162032412143e+17, 1.282162032512142e+17, 1.282162032612143e+17, 1.282162032712142e+17, 1.282162032812143e+17, 1.282162032912142e+17, 1.282162033012142e+17, 1.282162033112142e+17, 1.282162033212142e+17, 1.282162033312143e+17, 1.282162033412142e+17, 1.282162033512142e+17, 1.282162033612142e+17, 1.282162033712143e+17, 1.282162033812142e+17, 1.282162033912143e+17, 1.282162034012142e+17, 1.282162034112143e+17, 1.282162034212142e+17, 1.282162034312142e+17, 1.282162034412143e+17, 1.282162034512142e+17, 1.282162034612142e+17, 1.282162034712142e+17, 1.282162034812143e+17, 1.282162034912142e+17, 1.282162035012143e+17, 1.282162035112142e+17, 1.282162035212143e+17, 1.282162035312142e+17, 1.282162035412143e+17, 1.282162035512142e+17, 1.282162035612142e+17, 1.282162035712142e+17, 1.282162035812142e+17, 1.282162035912143e+17, 1.282162036012142e+17, 1.282162036112142e+17, 1.282162036212142e+17, 1.282162036312143e+17, 1.282162036412142e+17, 1.282162036512143e+17, 1.282162036612142e+17, 1.282162036712143e+17, 1.282162036812142e+17, 1.282162036912142e+17, 1.282162037012143e+17, 1.282162037112142e+17, 1.282162037212142e+17, 1.282162037312142e+17, 1.282162037412143e+17, 1.282162037512142e+17, 1.282162037612143e+17, 1.282162037712142e+17, 1.282162037812143e+17, 1.282162037912142e+17, 1.282162038012143e+17, 1.282162038112142e+17, 1.282162038212142e+17, 1.282162038312142e+17, 1.282162038412142e+17, 1.282162038512143e+17, 1.282162038612142e+17, 1.282162038712142e+17, 1.282162038812142e+17, 1.282162038912143e+17, 1.282162039012142e+17, 1.282162039112143e+17, 1.282162039212142e+17, 1.282162039312143e+17, 1.282162039412142e+17, 1.282162039512142e+17, 1.282162039612143e+17, 1.282162039712142e+17, 1.282162039812142e+17, 1.282162039912142e+17, 1.282162040012143e+17, 1.282162040112142e+17, 1.282162040212143e+17, 1.282162040312142e+17, 1.282162040412143e+17, 1.282162040512142e+17, 1.282162040612142e+17, 1.282162040712143e+17, 1.282162040812142e+17, 1.282162040912142e+17, 1.282162041012142e+17, 1.282162041112143e+17, 1.282162041212142e+17, 1.282162041312142e+17, 1.282162041412142e+17, 1.282162041512143e+17, 1.282162041612142e+17, 1.282162041712143e+17, 1.282162041812142e+17, 1.282162041912142e+17, 1.282162042012142e+17, 1.282162042112142e+17, 1.282162042212143e+17, 1.282162042312142e+17, 1.282162042412142e+17, 1.282162042512142e+17, 1.282162042612143e+17, 1.282162042712142e+17, 1.282162042812143e+17, 1.282162042912142e+17, 1.282162043012143e+17, 1.282162043112142e+17, 1.282162043212142e+17, 1.282162043312143e+17, 1.282162043412142e+17, 1.282162043512142e+17, 1.282162043612142e+17, 1.282162043712143e+17, 1.282162043812142e+17, 1.282162043912143e+17, 1.282162044012142e+17, 1.282162044112143e+17, 1.282162044212142e+17, 1.282162044312143e+17, 1.282162044412142e+17, 1.282162044512142e+17, 1.282162044612142e+17, 1.282162044712142e+17, 1.282162044812143e+17, 1.282162044912142e+17, 1.282162045012142e+17, 1.282162045112142e+17, 1.282162045212143e+17, 1.282162045312142e+17, 1.282162045412143e+17, 1.282162045512142e+17, 1.282162045612143e+17, 1.282162045712142e+17, 1.282162045812142e+17, 1.282162045912143e+17, 1.282162046012142e+17, 1.282162046112142e+17, 1.282162046212142e+17, 1.282162046312143e+17, 1.282162046412142e+17, 1.282162046512143e+17, 1.282162046612142e+17, 1.282162046712143e+17, 1.282162046812142e+17, 1.282162046912143e+17, 1.282162047012142e+17, 1.282162047112142e+17, 1.282162047212142e+17, 1.282162047312142e+17, 1.282162047412143e+17, 1.282162047512142e+17, 1.282162047612142e+17, 1.282162047712142e+17, 1.282162047812143e+17, 1.282162047912142e+17, 1.282162048012143e+17, 1.282162048112142e+17, 1.282162048212143e+17, 1.282162048312142e+17, 1.282162048412142e+17, 1.282162048512143e+17, 1.282162048612142e+17, 1.282162048712142e+17, 1.282162048812142e+17, 1.282162048912143e+17, 1.282162049012142e+17, 1.282162049112143e+17, 1.282162049212142e+17, 1.282162049312143e+17, 1.282162049412142e+17, 1.282162049512143e+17, 1.282162049612143e+17, 1.282162049712142e+17, 1.282162049812142e+17, 1.282162049912142e+17, 1.282162050012143e+17, 1.282162050112142e+17, 1.282162050212142e+17, 1.282162050312142e+17, 1.282162050412143e+17, 1.282162050512142e+17, 1.282162050612143e+17, 1.282162050712142e+17, 1.282162050812142e+17, 1.282162050912142e+17, 1.282162051012142e+17, 1.282162051112143e+17, 1.282162051212142e+17, 1.282162051312142e+17, 1.282162051412142e+17, 1.282162051512143e+17, 1.282162051612142e+17, 1.282162051712143e+17, 1.282162051812142e+17, 1.282162051912143e+17, 1.282162052012142e+17, 1.282162052112142e+17, 1.282162052212143e+17, 1.282162052312142e+17, 1.282162052412142e+17, 1.282162052512142e+17, 1.282162052612143e+17, 1.282162052712142e+17, 1.282162052812143e+17, 1.282162052912142e+17, 1.282162053012143e+17, 1.282162053112142e+17, 1.282162053212143e+17, 1.282162053312142e+17, 1.282162053412142e+17, 1.282162053512142e+17, 1.282162053612142e+17, 1.282162053712143e+17, 1.282162053812142e+17, 1.282162053912142e+17, 1.282162054012142e+17, 1.282162054112143e+17, 1.282162054212142e+17, 1.282162054312143e+17, 1.282162054412142e+17, 1.282162054512143e+17, 1.282162054612142e+17, 1.282162054712142e+17, 1.282162054812143e+17, 1.282162054912142e+17, 1.282162055012142e+17, 1.282162055112142e+17, 1.282162055212143e+17, 1.282162055312142e+17, 1.282162055412143e+17, 1.282162055512142e+17, 1.282162055612143e+17, 1.282162055712142e+17, 1.282162055812143e+17, 1.282162055912142e+17, 1.282162056012142e+17, 1.282162056112142e+17, 1.282162056212142e+17, 1.282162056312143e+17, 1.282162056412142e+17, 1.282162056512142e+17, 1.282162056612142e+17, 1.282162056712143e+17, 1.282162056812142e+17, 1.282162056912143e+17, 1.282162057012142e+17, 1.282162057112143e+17, 1.282162057212142e+17, 1.282162057312142e+17, 1.282162057412143e+17, 1.282162057512142e+17, 1.282162057612142e+17, 1.282162057712142e+17, 1.282162057812143e+17, 1.282162057912142e+17, 1.282162058012143e+17, 1.282162058112142e+17, 1.282162058212143e+17, 1.282162058312142e+17, 1.282162058412143e+17, 1.282162058512142e+17, 1.282162058612142e+17, 1.282162058712142e+17, 1.282162058812142e+17, 1.282162058912143e+17, 1.282162059012142e+17, 1.282162059112142e+17, 1.282162059212142e+17, 1.282162059312143e+17, 1.282162059412142e+17, 1.282162059512143e+17, 1.282162059612142e+17, 1.282162059712143e+17, 1.282162059812142e+17, 1.282162059912142e+17, 1.282162060012143e+17, 1.282162060112142e+17, 1.282162060212142e+17, 1.282162060312142e+17, 1.282162060412143e+17, 1.282162060512142e+17, 1.282162060612143e+17, 1.282162060712142e+17, 1.282162060812143e+17, 1.282162060912142e+17, 1.282162061012142e+17, 1.282162061112143e+17, 1.282162061212142e+17, 1.282162061312142e+17, 1.282162061412142e+17, 1.282162061512143e+17, 1.282162061612142e+17, 1.282162061712143e+17, 1.282162061812142e+17, 1.282162061912143e+17, 1.282162062012142e+17, 1.282162062112143e+17, 1.282162062212142e+17, 1.282162062312142e+17, 1.282162062412142e+17, 1.282162062512142e+17, 1.282162062612143e+17, 1.282162062712142e+17, 1.282162062812142e+17, 1.282162062912142e+17, 1.282162063012143e+17, 1.282162063112142e+17, 1.282162063212143e+17, 1.282162063312142e+17, 1.282162063412143e+17, 1.282162063512142e+17, 1.282162063612142e+17, 1.282162063712143e+17, 1.282162063812142e+17, 1.282162063912142e+17, 1.282162064012142e+17, 1.282162064112143e+17, 1.282162064212142e+17, 1.282162064312143e+17, 1.282162064412142e+17, 1.282162064512143e+17, 1.282162064612142e+17, 1.282162064712143e+17, 1.282162064812142e+17, 1.282162064912142e+17, 1.282162065012142e+17, 1.282162065112142e+17, 1.282162065212143e+17, 1.282162065312142e+17, 1.282162065412142e+17, 1.282162065512142e+17, 1.282162065612143e+17, 1.282162065712142e+17, 1.282162065812143e+17, 1.282162065912142e+17, 1.282162066012143e+17, 1.282162066112142e+17, 1.282162066212142e+17, 1.282162066312143e+17, 1.282162066412142e+17, 1.282162066512142e+17, 1.282162066612142e+17, 1.282162066712143e+17, 1.282162066812142e+17, 1.282162066912143e+17, 1.282162067012142e+17, 1.282162067112143e+17, 1.282162067212142e+17, 1.282162067312143e+17, 1.282162067412142e+17, 1.282162067512142e+17, 1.282162067612142e+17, 1.282162067712142e+17, 1.282162067812143e+17, 1.282162067912142e+17, 1.282162068012142e+17, 1.282162068112142e+17, 1.282162068212143e+17, 1.282162068312142e+17, 1.282162068412143e+17, 1.282162068512142e+17, 1.282162068612143e+17, 1.282162068712142e+17, 1.282162068812142e+17, 1.282162068912143e+17, 1.282162069012142e+17, 1.282162069112142e+17, 1.282162069212142e+17, 1.282162069312143e+17, 1.282162069412142e+17, 1.282162069512143e+17, 1.282162069612142e+17, 1.282162069712143e+17, 1.282162069812142e+17, 1.282162069912142e+17, 1.282162070012143e+17, 1.282162070112142e+17, 1.282162070212142e+17, 1.282162070312142e+17, 1.282162070412143e+17, 1.282162070512142e+17, 1.282162070612142e+17, 1.282162070712142e+17, 1.282162070812143e+17, 1.282162070912142e+17, 1.282162071012143e+17, 1.282162071112142e+17, 1.282162071212142e+17, 1.282162071312142e+17, 1.282162071412142e+17, 1.282162071512143e+17, 1.282162071612142e+17, 1.282162071712142e+17, 1.282162071812142e+17, 1.282162071912143e+17, 1.282162072012142e+17, 1.282162072112143e+17, 1.282162072212142e+17, 1.282162072312143e+17, 1.282162072412142e+17, 1.282162072512142e+17, 1.282162072612143e+17, 1.282162072712142e+17, 1.282162072812142e+17, 1.282162072912142e+17, 1.282162073012143e+17, 1.282162073112142e+17, 1.282162073212143e+17, 1.282162073312142e+17, 1.282162073412143e+17, 1.282162073512142e+17, 1.282162073612143e+17, 1.282162073712142e+17, 1.282162073812142e+17, 1.282162073912142e+17, 1.282162074012142e+17, 1.282162074112143e+17, 1.282162074212142e+17, 1.282162074312142e+17, 1.282162074412142e+17, 1.282162074512143e+17, 1.282162074612142e+17, 1.282162074712143e+17, 1.282162074812142e+17, 1.282162074912143e+17, 1.282162075012142e+17, 1.282162075112142e+17, 1.282162075212143e+17, 1.282162075312142e+17, 1.282162075412142e+17, 1.282162075512142e+17, 1.282162075612143e+17, 1.282162075712142e+17, 1.282162075812143e+17, 1.282162075912142e+17, 1.282162076012143e+17, 1.282162076112142e+17, 1.282162076212143e+17, 1.282162076312142e+17, 1.282162076412142e+17, 1.282162076512142e+17, 1.282162076612142e+17, 1.282162076712143e+17, 1.282162076812142e+17, 1.282162076912142e+17, 1.282162077012142e+17, 1.282162077112143e+17, 1.282162077212142e+17, 1.282162077312143e+17, 1.282162077412142e+17, 1.282162077512143e+17, 1.282162077612142e+17, 1.282162077712142e+17, 1.282162077812143e+17, 1.282162077912142e+17, 1.282162078012142e+17, 1.282162078112142e+17, 1.282162078212143e+17, 1.282162078312142e+17, 1.282162078412143e+17, 1.282162078512142e+17, 1.282162078612143e+17, 1.282162078712142e+17, 1.282162078812143e+17, 1.282162078912143e+17, 1.282162079012142e+17, 1.282162079112142e+17, 1.282162079212142e+17, 1.282162079312143e+17, 1.282162079412142e+17, 1.282162079512142e+17, 1.282162079612142e+17, 1.282162079712143e+17, 1.282162079812142e+17, 1.282162079912143e+17, 1.282162080012142e+17, 1.282162080112142e+17, 1.282162080212142e+17, 1.282162080312142e+17, 1.282162080412143e+17, 1.282162080512142e+17, 1.282162080612142e+17, 1.282162080712142e+17, 1.282162080812143e+17, 1.282162080912142e+17, 1.282162081012143e+17, 1.282162081112142e+17, 1.282162081212143e+17, 1.282162081312142e+17, 1.282162081412142e+17, 1.282162081512143e+17, 1.282162081612142e+17, 1.282162081712142e+17, 1.282162081812142e+17, 1.282162081912143e+17, 1.282162082012142e+17, 1.282162082112143e+17, 1.282162082212142e+17, 1.282162082312143e+17, 1.282162082412142e+17, 1.282162082512143e+17, 1.282162082612142e+17, 1.282162082712142e+17, 1.282162082812142e+17, 1.282162082912142e+17, 1.282162083012143e+17, 1.282162083112142e+17, 1.282162083212142e+17, 1.282162083312142e+17, 1.282162083412143e+17, 1.282162083512142e+17, 1.282162083612143e+17, 1.282162083712142e+17, 1.282162083812143e+17, 1.282162083912142e+17, 1.282162084012142e+17, 1.282162084112143e+17, 1.282162084212142e+17, 1.282162084312142e+17, 1.282162084412142e+17, 1.282162084512143e+17, 1.282162084612142e+17, 1.282162084712143e+17, 1.282162084812142e+17, 1.282162084912143e+17, 1.282162085012142e+17, 1.282162085112143e+17, 1.282162085212142e+17, 1.282162085312142e+17, 1.282162085412142e+17, 1.282162085512142e+17, 1.282162085612143e+17, 1.282162085712142e+17, 1.282162085812142e+17, 1.282162085912142e+17, 1.282162086012143e+17, 1.282162086112142e+17, 1.282162086212143e+17, 1.282162086312142e+17, 1.282162086412143e+17, 1.282162086512142e+17, 1.282162086612142e+17, 1.282162086712143e+17, 1.282162086812142e+17, 1.282162086912142e+17, 1.282162087012142e+17, 1.282162087112143e+17, 1.282162087212142e+17, 1.282162087312143e+17, 1.282162087412142e+17, 1.282162087512143e+17, 1.282162087612142e+17, 1.282162087712143e+17, 1.282162087812142e+17, 1.282162087912142e+17, 1.282162088012142e+17, 1.282162088112142e+17, 1.282162088212143e+17, 1.282162088312142e+17, 1.282162088412142e+17, 1.282162088512142e+17, 1.282162088612143e+17, 1.282162088712142e+17, 1.282162088812143e+17, 1.282162088912142e+17, 1.282162089012142e+17, 1.282162089112142e+17, 1.282162089212142e+17, 1.282162089312143e+17, 1.282162089412142e+17, 1.282162089512142e+17, 1.282162089612142e+17, 1.282162089712143e+17, 1.282162089812142e+17, 1.282162089912143e+17, 1.282162090012142e+17, 1.282162090112143e+17, 1.282162090212142e+17, 1.282162090312142e+17, 1.282162090412143e+17, 1.282162090512142e+17, 1.282162090612142e+17, 1.282162090712142e+17, 1.282162090812143e+17, 1.282162090912142e+17, 1.282162091012143e+17, 1.282162091112142e+17, 1.282162091212143e+17, 1.282162091312142e+17, 1.282162091412143e+17, 1.282162091512142e+17, 1.282162091612142e+17, 1.282162091712142e+17, 1.282162091812142e+17, 1.282162091912143e+17, 1.282162092012142e+17, 1.282162092112142e+17, 1.282162092212142e+17, 1.282162092312143e+17, 1.282162092412142e+17, 1.282162092512143e+17, 1.282162092612142e+17, 1.282162092712143e+17, 1.282162092812142e+17, 1.282162092912142e+17, 1.282162093012143e+17, 1.282162093112142e+17, 1.282162093212142e+17, 1.282162093312142e+17, 1.282162093412143e+17, 1.282162093512142e+17, 1.282162093612143e+17, 1.282162093712142e+17, 1.282162093812143e+17, 1.282162093912142e+17, 1.282162094012143e+17, 1.282162094112142e+17, 1.282162094212142e+17, 1.282162094312142e+17, 1.282162094412142e+17, 1.282162094512143e+17, 1.282162094612142e+17, 1.282162094712142e+17, 1.282162094812142e+17, 1.282162094912143e+17, 1.282162095012142e+17, 1.282162095112143e+17, 1.282162095212142e+17, 1.282162095312143e+17, 1.282162095412142e+17, 1.282162095512142e+17, 1.282162095612143e+17, 1.282162095712142e+17, 1.282162095812142e+17, 1.282162095912142e+17, 1.282162096012143e+17, 1.282162096112142e+17, 1.282162096212143e+17, 1.282162096312142e+17, 1.282162096412143e+17, 1.282162096512142e+17, 1.282162096612143e+17, 1.282162096712142e+17, 1.282162096812142e+17, 1.282162096912142e+17, 1.282162097012142e+17, 1.282162097112143e+17, 1.282162097212142e+17, 1.282162097312142e+17, 1.282162097412142e+17, 1.282162097512143e+17, 1.282162097612142e+17, 1.282162097712143e+17, 1.282162097812142e+17, 1.282162097912143e+17, 1.282162098012142e+17, 1.282162098112142e+17, 1.282162098212143e+17, 1.282162098312142e+17, 1.282162098412142e+17, 1.282162098512142e+17, 1.282162098612143e+17, 1.282162098712142e+17, 1.282162098812143e+17, 1.282162098912142e+17, 1.282162099012143e+17, 1.282162099112142e+17, 1.282162099212142e+17, 1.282162099312143e+17, 1.282162099412142e+17, 1.282162099512142e+17, 1.282162099612142e+17, 1.282162099712143e+17, 1.282162099812142e+17, 1.282162099912143e+17, 1.282162100012142e+17, 1.282162100112143e+17, 1.282162100212142e+17, 1.282162100312143e+17, 1.282162100412142e+17, 1.282162100512142e+17, 1.282162100612142e+17, 1.282162100712142e+17, 1.282162100812143e+17, 1.282162100912142e+17, 1.282162101012142e+17, 1.282162101112142e+17, 1.282162101212143e+17, 1.282162101312142e+17, 1.282162101412143e+17, 1.282162101512142e+17, 1.282162101612143e+17, 1.282162101712142e+17, 1.282162101812142e+17, 1.282162101912143e+17, 1.282162102012142e+17, 1.282162102112142e+17, 1.282162102212142e+17, 1.282162102312143e+17, 1.282162102412142e+17, 1.282162102512143e+17, 1.282162102612142e+17, 1.282162102712143e+17, 1.282162102812142e+17, 1.282162102912143e+17, 1.282162103012142e+17, 1.282162103112142e+17, 1.282162103212142e+17, 1.282162103312142e+17, 1.282162103412143e+17, 1.282162103512142e+17, 1.282162103612142e+17, 1.282162103712142e+17, 1.282162103812143e+17, 1.282162103912142e+17, 1.282162104012143e+17, 1.282162104112142e+17, 1.282162104212143e+17, 1.282162104312142e+17, 1.282162104412142e+17, 1.282162104512143e+17, 1.282162104612142e+17, 1.282162104712142e+17, 1.282162104812142e+17, 1.282162104912143e+17, 1.282162105012142e+17, 1.282162105112143e+17, 1.282162105212142e+17, 1.282162105312143e+17, 1.282162105412142e+17, 1.282162105512143e+17, 1.282162105612142e+17, 1.282162105712142e+17, 1.282162105812142e+17, 1.282162105912142e+17, 1.282162106012143e+17, 1.282162106112142e+17, 1.282162106212142e+17, 1.282162106312142e+17, 1.282162106412143e+17, 1.282162106512142e+17, 1.282162106612143e+17, 1.282162106712142e+17, 1.282162106812143e+17, 1.282162106912142e+17, 1.282162107012142e+17, 1.282162107112143e+17, 1.282162107212142e+17, 1.282162107312142e+17, 1.282162107412142e+17, 1.282162107512143e+17, 1.282162107612142e+17, 1.282162107712143e+17, 1.282162107812142e+17, 1.282162107912143e+17, 1.282162108012142e+17, 1.282162108112142e+17, 1.282162108212143e+17, 1.282162108312142e+17, 1.282162108412142e+17, 1.282162108512142e+17, 1.282162108612143e+17, 1.282162108712142e+17, 1.282162108812142e+17, 1.282162108912142e+17, 1.282162109012143e+17, 1.282162109112142e+17, 1.282162109212143e+17, 1.282162109312142e+17, 1.282162109412142e+17, 1.282162109512142e+17, 1.282162109612142e+17, 1.282162109712143e+17, 1.282162109812142e+17, 1.282162109912142e+17, 1.282162110012142e+17, 1.282162110112143e+17, 1.282162110212142e+17, 1.282162110312143e+17, 1.282162110412142e+17, 1.282162110512143e+17, 1.282162110612142e+17, 1.282162110712142e+17, 1.282162110812143e+17, 1.282162110912142e+17, 1.282162111012142e+17, 1.282162111112142e+17, 1.282162111212143e+17, 1.282162111312142e+17, 1.282162111412143e+17, 1.282162111512142e+17, 1.282162111612143e+17, 1.282162111712142e+17, 1.282162111812143e+17, 1.282162111912142e+17, 1.282162112012142e+17, 1.282162112112142e+17, 1.282162112212142e+17, 1.282162112312143e+17, 1.282162112412142e+17, 1.282162112512142e+17, 1.282162112612142e+17, 1.282162112712143e+17, 1.282162112812142e+17, 1.282162112912143e+17, 1.282162113012142e+17, 1.282162113112143e+17, 1.282162113212142e+17, 1.282162113312142e+17, 1.282162113412143e+17, 1.282162113512142e+17, 1.282162113612142e+17, 1.282162113712142e+17, 1.282162113812143e+17, 1.282162113912142e+17, 1.282162114012143e+17, 1.282162114112142e+17, 1.282162114212143e+17, 1.282162114312142e+17, 1.282162114412143e+17, 1.282162114512142e+17, 1.282162114612142e+17, 1.282162114712142e+17, 1.282162114812142e+17, 1.282162114912143e+17, 1.282162115012142e+17, 1.282162115112142e+17, 1.282162115212142e+17, 1.282162115312143e+17, 1.282162115412142e+17, 1.282162115512143e+17, 1.282162115612142e+17, 1.282162115712143e+17, 1.282162115812142e+17, 1.282162115912142e+17, 1.282162116012143e+17, 1.282162116112142e+17, 1.282162116212142e+17, 1.282162116312142e+17, 1.282162116412143e+17, 1.282162116512142e+17, 1.282162116612143e+17, 1.282162116712142e+17, 1.282162116812143e+17, 1.282162116912142e+17, 1.282162117012143e+17, 1.282162117112143e+17, 1.282162117212142e+17, 1.282162117312142e+17, 1.282162117412142e+17, 1.282162117512143e+17, 1.282162117612142e+17, 1.282162117712142e+17, 1.282162117812142e+17, 1.282162117912143e+17, 1.282162118012142e+17, 1.282162118112143e+17, 1.282162118212142e+17, 1.282162118312142e+17, 1.282162118412142e+17, 1.282162118512142e+17, 1.282162118612143e+17, 1.282162118712142e+17, 1.282162118812142e+17, 1.282162118912142e+17, 1.282162119012143e+17, 1.282162119112142e+17, 1.282162119212143e+17, 1.282162119312142e+17, 1.282162119412143e+17, 1.282162119512142e+17, 1.282162119612142e+17, 1.282162119712143e+17, 1.282162119812142e+17, 1.282162119912142e+17, 1.282162120012142e+17, 1.282162120112143e+17, 1.282162120212142e+17, 1.282162120312143e+17, 1.282162120412142e+17, 1.282162120512143e+17, 1.282162120612142e+17, 1.282162120712143e+17, 1.282162120812142e+17, 1.282162120912142e+17, 1.282162121012142e+17},
			             {1.282162157812142e+17, 1.282162157912143e+17, 1.282162158012142e+17, 1.282162158112142e+17, 1.282162158212142e+17};
			mask_depths = {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}, {}}, {{}, {}, {}, {}, {}};
		}
	}
}
