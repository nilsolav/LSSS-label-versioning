netcdf mask {
	:date_created = "20200811T114628";
	:mask_convention_version = "0.1";
	:mask_convention_name = "SONAR-netCDF4";
	:mask_convention_authority = "ICES, IMR";
	:rights = "Unrestricted rights";
	:license = "None";
	:Conventions = "CF-1.7, ACDD-1.3, SONAR-netCDF4-2.0";
	:keywords = "scrutinisation mask, echosounder";
	:summary = "Contains definitions of echogram scrutiny masks";
	:title = "Echogram scrutiny masks";

group: Interpretation {
	group: v1{
		:version = "1";
		:version_save_date = "20200811T114628";
		:version_author = "GJM";
		:version_comment = "Initial scrutiny";
		types:
			byte enum region_t {empty_water = 0, no_data = 1, analysis = 2, track = 3, marker = 4};
			byte enum region_dim_t {twoD = 0, threeD = 1};
			float(*) mask_depth_t;
			mask_depth_t(*) mask_depths_t;
			uint64(*) mask_time_t;
		dimensions:
			regions = 1;
			channels = 4;
			categories = 4;
		variables:
			float sound_speed;
				sound_speed:long_name = "Sound speed used to convert echo time into range";
				sound_speed:standard_name = "speed_of_sound_in_sea_water";
				sound_speed:units = "m/s";
				sound_speed:valid_min = 0.0f;

			// The bounding box of each region
			float min_depth(regions);
				min_depth:long_name = "Minimum depth for each region";
				min_depth:units = "m";
				min_depth:valid_min = 0.0f;
			float max_depth(regions);
				max_depth:long_name = "Maximum depth for each regions";
				max_depth:units = "m";
				max_depth:valid_min = 0.0f;
			uint64 start_time(regions);
				start_time:long_name = "Timestamp of the earliest data point in each region";
				start_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				start_time:axis = "T";
				start_time:calendar = "gregorian";
				start_time:standard_name = "time";
			uint64 end_time(regions);
				end_time:long_name = "Timestamp of the latest data point in each region";
				end_time:units = "milliseconds since 1601-01-01 00:00:00Z";
				end_time:axis = "T";
				end_time:calendar = "gregorian";
				end_time:standard_name = "time";
				
			region_dim_t region_dimension; 
				region_dimension:long_name = "Region dimension";

			int region_id(regions);
				region_id:long_name = "Dataset-unique identification number for each region";
			string region_name(regions);
				region_name:long_name = "Name of each region";
				region_name:_Encoding = "utf-8";
			string region_provenance(regions);
				region_provenance:long_name = "Provenance of each region"; 
				region_provenance:_Encoding = "utf-8";
			string region_comment(regions);
				region_comment:long_name = "Comment for each region";
				region_comment:_Encoding = "utf-8";
			int region_order(regions);
				region_order:long_name = "The stacking order of the region";
				region_order:comment = "Regions of the same order cannot overlap";
			region_t region_type(regions);
				region_type:long_name = "Region type";
			
			// The acosutic categories. Each layer may have several categories and proportions.
			string region_category_names(categories);
				region_category_names:long_name = "Categorisation name";
				region_category_names:_Encoding = "utf-8";
			float region_category_proportions(categories);
				region_category_proportions:long_name = "Proportion of backscatter for the categorisation";
				region_category_proportions:value_range = 0.0f, 1.0f;
			int region_category_ids(categories);
				region_category_ids:long_name = "region_id of this categorisation and proportion";
			
			string channel_names(channels);
				channel_names:long_name = "Echosounder channel names";
				channel_names:_Encoding = "utf-8";
			uint region_channels(regions);
				region_channels:long_name = "Echosounder channels that this region applies to";
				region_channels:description = "Bit mask derived from channel_names (index 1 of channel_names = bit 1, index 2 = bit 2, etc). Set bits in excess of the number of channels are to be ignored.";
				region_channels:_FillValue = 4294967295; // 2^32-1
				
			mask_time_t mask_times(regions);
				mask_times:long_name = "Timestamp of each mask point";
				mask_times:units = "milliseconds since 1601-01-01 00:00:00Z";
				mask_times:axis = "T";
				mask_times:calendar = "gregorian";
				mask_times:standard_name = "time";
			mask_depths_t mask_depths(regions);
				mask_depths:long_name = "Depth pairs of mask";
				mask_depths:units = "m";
				mask_depths:valid_min = 0.0f;

		data:
			region_dimension = twoD;
			sound_speed = 1496;
			min_depth =  46.8;
			max_depth =  54.6;
			start_time = 129162944163945344;
			end_time = 129162944276601600;
			region_id = 1;
			region_name = "Layer1";
			region_provenance = "LSSS";
			region_comment = "";
			region_category_names = "1", "1", "1", "1";
			region_category_proportions = 1.0, 1.0, 1.0, 1.0;
			region_category_ids = 1, 2, 3, 4;
			region_type = analysis;
			channel_names = "18", "38", "120", "200";
			region_channels = 15;
			mask_times = {1.291629441639453e+17, 1.291629441672266e+17, 1.291629441703516e+17, 1.291629441736329e+17, 1.29162944176914e+17, 1.291629441800392e+17, 1.291629441833203e+17, 1.291629441864453e+17, 1.291629441897266e+17, 1.291629441928516e+17, 1.291629441961329e+17, 1.29162944199414e+17, 1.291629442025391e+17, 1.291629442058204e+17, 1.291629442089453e+17, 1.291629442122266e+17, 1.291629442155078e+17, 1.291629442186328e+17, 1.291629442219141e+17, 1.291629442250391e+17, 1.291629442283204e+17, 1.291629442316015e+17, 1.291629442347267e+17, 1.291629442380079e+17, 1.291629442411328e+17, 1.291629442444141e+17, 1.291629442476954e+17, 1.291629442508204e+17, 1.291629442541015e+17, 1.291629442572266e+17, 1.291629442605079e+17, 1.291629442636328e+17, 1.29162944266914e+17, 1.291629442701953e+17, 1.291629442733203e+17, 1.291629442766016e+17};
			mask_depths = {{51.6, 54.6}, {51.6, 54.6}, {51.6, 54.6}, {51.5, 51.6, 54.6}, {51.2, 51.4, 54.6}, {51.1, 51.2, 54.6}, {50.2, 50.9, 54.6}, {49.4, 50.0, 54.6}, {49.0, 49.3, 54.6}, {48.5, 48.9, 54.5}, {47.9, 48.5, 54.5}, {47.7, 54.5}, {47.6, 54.5}, {47.5, 54.5}, {47.4, 54.5}, {47.3, 54.5}, {47.2, 54.6}, {47.1, 54.6}, {47.0, 54.6}, {46.8, 54.6}, {46.8, 54.6}, {46.8, 54.6}, {46.9, 54.6}, {46.8, 46.9, 54.6}, {46.8, 54.6}, {46.9, 47.0, 54.6}, {47.2, 47.4, 54.6}, {47.6, 47.9, 54.6}, {48.1, 54.6}, {48.6, 54.6}, {48.7, 54.6}, {48.8, 54.6}, {48.9, 49.1, 54.5}, {49.5, 50.2, 54.5}, {50.4, 52.5, 54.5}, {52.5, 54.5}};
		}
	}
}
